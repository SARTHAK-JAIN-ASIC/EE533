module weight_rom (
    input clk,
    input reset,
    output [15:0] data_out_0,
	output [15:0] data_out_1,
	output [15:0] data_out_2,
	output [15:0] data_out_3,
	output [15:0] data_out_4,
	output [15:0] data_out_5,
	output [15:0] data_out_6,
	output [15:0] data_out_7,
	output [15:0] data_out_8,
	output [15:0] data_out_9,
	output [15:0] data_out_10,
	output [15:0] data_out_11,
	output [15:0] data_out_12,
	output [15:0] data_out_13,
	output [15:0] data_out_14,
	output [15:0] data_out_15,
	output [15:0] data_out_16,
	output [15:0] data_out_17,
	output [15:0] data_out_18,
	output [15:0] data_out_19,
	output [15:0] data_out_20,
	output [15:0] data_out_21,
	output [15:0] data_out_22,
	output [15:0] data_out_23,
	output [15:0] data_out_24,
	output [15:0] data_out_25,
	output [15:0] data_out_26,
	output [15:0] data_out_27,
	output [15:0] data_out_28,
	output [15:0] data_out_29,
	output [15:0] data_out_30,
	output [15:0] data_out_31,
	output [15:0] data_out_32,
	output [15:0] data_out_33,
	output [15:0] data_out_34,
	output [15:0] data_out_35,
	output [15:0] data_out_36,
	output [15:0] data_out_37,
	output [15:0] data_out_38,
	output [15:0] data_out_39,
	output [15:0] data_out_40,
	output [15:0] data_out_41,
	output [15:0] data_out_42,
	output [15:0] data_out_43,
	output [15:0] data_out_44,
	output [15:0] data_out_45,
	output [15:0] data_out_46,
	output [15:0] data_out_47,
	output [15:0] data_out_48,
	output [15:0] data_out_49,
	output [15:0] data_out_50,
	output [15:0] data_out_51,
	output [15:0] data_out_52,
	output [15:0] data_out_53,
	output [15:0] data_out_54,
	output [15:0] data_out_55,
	output [15:0] data_out_56,
	output [15:0] data_out_57,
	output [15:0] data_out_58,
	output [15:0] data_out_59,
	output [15:0] data_out_60,
	output [15:0] data_out_61,
	output [15:0] data_out_62,
	output [15:0] data_out_63,
	output [15:0] data_out_64,
	output [15:0] data_out_65,
	output [15:0] data_out_66,
	output [15:0] data_out_67,
	output [15:0] data_out_68,
	output [15:0] data_out_69,
	output [15:0] data_out_70,
	output [15:0] data_out_71,
	output [15:0] data_out_72,
	output [15:0] data_out_73,
	output [15:0] data_out_74,
	output [15:0] data_out_75,
	output [15:0] data_out_76,
	output [15:0] data_out_77,
	output [15:0] data_out_78,
	output [15:0] data_out_79,
	output [15:0] data_out_80,
	output [15:0] data_out_81,
	output [15:0] data_out_82,
	output [15:0] data_out_83,
	output [15:0] data_out_84,
	output [15:0] data_out_85,
	output [15:0] data_out_86,
	output [15:0] data_out_87,
	output [15:0] data_out_88,
	output [15:0] data_out_89,
	output [15:0] data_out_90,
	output [15:0] data_out_91,
	output [15:0] data_out_92,
	output [15:0] data_out_93,
	output [15:0] data_out_94,
	output [15:0] data_out_95,
	output [15:0] data_out_96,
	output [15:0] data_out_97,
	output [15:0] data_out_98,
	output [15:0] data_out_99,
	output [15:0] data_out_100,
	output [15:0] data_out_101,
	output [15:0] data_out_102,
	output [15:0] data_out_103,
	output [15:0] data_out_104,
	output [15:0] data_out_105,
	output [15:0] data_out_106,
	output [15:0] data_out_107,
	output [15:0] data_out_108,
	output [15:0] data_out_109,
	output [15:0] data_out_110,
	output [15:0] data_out_111,
	output [15:0] data_out_112,
	output [15:0] data_out_113,
	output [15:0] data_out_114,
	output [15:0] data_out_115,
	output [15:0] data_out_116,
	output [15:0] data_out_117,
	output [15:0] data_out_118,
	output [15:0] data_out_119,
	output [15:0] data_out_120,
	output [15:0] data_out_121,
	output [15:0] data_out_122,
	output [15:0] data_out_123,
	output [15:0] data_out_124,
	output [15:0] data_out_125,
	output [15:0] data_out_126,
	output [15:0] data_out_127,
	output [15:0] data_out_128,
	output [15:0] data_out_129,
	output [15:0] data_out_130,
	output [15:0] data_out_131,
	output [15:0] data_out_132,
	output [15:0] data_out_133,
	output [15:0] data_out_134,
	output [15:0] data_out_135,
	output [15:0] data_out_136,
	output [15:0] data_out_137,
	output [15:0] data_out_138,
	output [15:0] data_out_139,
	output [15:0] data_out_140,
	output [15:0] data_out_141,
	output [15:0] data_out_142,
	output [15:0] data_out_143,
	output [15:0] data_out_144,
	output [15:0] data_out_145,
	output [15:0] data_out_146,
	output [15:0] data_out_147,
	output [15:0] data_out_148,
	output [15:0] data_out_149,
	output [15:0] data_out_150,
	output [15:0] data_out_151,
	output [15:0] data_out_152,
	output [15:0] data_out_153,
	output [15:0] data_out_154,
	output [15:0] data_out_155,
	output [15:0] data_out_156,
	output [15:0] data_out_157,
	output [15:0] data_out_158,
	output [15:0] data_out_159,
	output [15:0] data_out_160,
	output [15:0] data_out_161,
	output [15:0] data_out_162,
	output [15:0] data_out_163,
	output [15:0] data_out_164,
	output [15:0] data_out_165,
	output [15:0] data_out_166,
	output [15:0] data_out_167,
	output [15:0] data_out_168,
	output [15:0] data_out_169,
	output [15:0] data_out_170,
	output [15:0] data_out_171,
	output [15:0] data_out_172,
	output [15:0] data_out_173,
	output [15:0] data_out_174,
	output [15:0] data_out_175,
	output [15:0] data_out_176,
	output [15:0] data_out_177,
	output [15:0] data_out_178,
	output [15:0] data_out_179,
	output [15:0] data_out_180,
	output [15:0] data_out_181,
	output [15:0] data_out_182,
	output [15:0] data_out_183,
	output [15:0] data_out_184,
	output [15:0] data_out_185,
	output [15:0] data_out_186,
	output [15:0] data_out_187,
	output [15:0] data_out_188,
	output [15:0] data_out_189,
	output [15:0] data_out_190,
	output [15:0] data_out_191,
	output [15:0] data_out_192,
	output [15:0] data_out_193,
	output [15:0] data_out_194,
	output [15:0] data_out_195,
	output [15:0] data_out_196,
	output [15:0] data_out_197,
	output [15:0] data_out_198,
	output [15:0] data_out_199,
	output [15:0] data_out_200,
	output [15:0] data_out_201,
	output [15:0] data_out_202,
	output [15:0] data_out_203,
	output [15:0] data_out_204,
	output [15:0] data_out_205,
	output [15:0] data_out_206,
	output [15:0] data_out_207,
	output [15:0] data_out_208,
	output [15:0] data_out_209,
	output [15:0] data_out_210,
	output [15:0] data_out_211,
	output [15:0] data_out_212,
	output [15:0] data_out_213,
	output [15:0] data_out_214,
	output [15:0] data_out_215,
	output [15:0] data_out_216,
	output [15:0] data_out_217,
	output [15:0] data_out_218,
	output [15:0] data_out_219,
	output [15:0] data_out_220,
	output [15:0] data_out_221,
	output [15:0] data_out_222,
	output [15:0] data_out_223,
	output [15:0] data_out_224,
	output [15:0] data_out_225,
	output [15:0] data_out_226,
	output [15:0] data_out_227,
	output [15:0] data_out_228,
	output [15:0] data_out_229,
	output [15:0] data_out_230,
	output [15:0] data_out_231,
	output [15:0] data_out_232,
	output [15:0] data_out_233,
	output [15:0] data_out_234,
	output [15:0] data_out_235,
	output [15:0] data_out_236,
	output [15:0] data_out_237,
	output [15:0] data_out_238,
	output [15:0] data_out_239,
	output [15:0] data_out_240,
	output [15:0] data_out_241,
	output [15:0] data_out_242,
	output [15:0] data_out_243,
	output [15:0] data_out_244,
	output [15:0] data_out_245,
	output [15:0] data_out_246,
	output [15:0] data_out_247,
	output [15:0] data_out_248,
	output [15:0] data_out_249,
	output [15:0] data_out_250,
	output [15:0] data_out_251,
	output [15:0] data_out_252,
	output [15:0] data_out_253,
	output [15:0] data_out_254,
	output [15:0] data_out_255,
	output [15:0] data_out_256,
	output [15:0] data_out_257,
	output [15:0] data_out_258,
	output [15:0] data_out_259,
	output [15:0] data_out_260,
	output [15:0] data_out_261,
	output [15:0] data_out_262,
	output [15:0] data_out_263,
	output [15:0] data_out_264,
	output [15:0] data_out_265,
	output [15:0] data_out_266,
	output [15:0] data_out_267,
	output [15:0] data_out_268,
	output [15:0] data_out_269,
	output [15:0] data_out_270,
	output [15:0] data_out_271,
	output [15:0] data_out_272,
	output [15:0] data_out_273,
	output [15:0] data_out_274,
	output [15:0] data_out_275,
	output [15:0] data_out_276,
	output [15:0] data_out_277,
	output [15:0] data_out_278,
	output [15:0] data_out_279,
	output [15:0] data_out_280,
	output [15:0] data_out_281,
	output [15:0] data_out_282,
	output [15:0] data_out_283,
	output [15:0] data_out_284,
	output [15:0] data_out_285,
	output [15:0] data_out_286,
	output [15:0] data_out_287,
	output [15:0] data_out_288,
	output [15:0] data_out_289,
	output [15:0] data_out_290,
	output [15:0] data_out_291,
	output [15:0] data_out_292,
	output [15:0] data_out_293,
	output [15:0] data_out_294,
	output [15:0] data_out_295,
	output [15:0] data_out_296,
	output [15:0] data_out_297,
	output [15:0] data_out_298,
	output [15:0] data_out_299,
	output [15:0] data_out_300,
	output [15:0] data_out_301,
	output [15:0] data_out_302,
	output [15:0] data_out_303,
	output [15:0] data_out_304,
	output [15:0] data_out_305,
	output [15:0] data_out_306,
	output [15:0] data_out_307,
	output [15:0] data_out_308,
	output [15:0] data_out_309,
	output [15:0] data_out_310,
	output [15:0] data_out_311,
	output [15:0] data_out_312,
	output [15:0] data_out_313,
	output [15:0] data_out_314,
	output [15:0] data_out_315,
	output [15:0] data_out_316,
	output [15:0] data_out_317,
	output [15:0] data_out_318,
	output [15:0] data_out_319,
	output [15:0] data_out_320,
	output [15:0] data_out_321,
	output [15:0] data_out_322,
	output [15:0] data_out_323,
	output [15:0] data_out_324,
	output [15:0] data_out_325,
	output [15:0] data_out_326,
	output [15:0] data_out_327,
	output [15:0] data_out_328,
	output [15:0] data_out_329,
	output [15:0] data_out_330,
	output [15:0] data_out_331,
	output [15:0] data_out_332,
	output [15:0] data_out_333,
	output [15:0] data_out_334,
	output [15:0] data_out_335,
	output [15:0] data_out_336,
	output [15:0] data_out_337,
	output [15:0] data_out_338,
	output [15:0] data_out_339,
	output [15:0] data_out_340,
	output [15:0] data_out_341,
	output [15:0] data_out_342,
	output [15:0] data_out_343,
	output [15:0] data_out_344,
	output [15:0] data_out_345,
	output [15:0] data_out_346,
	output [15:0] data_out_347,
	output [15:0] data_out_348,
	output [15:0] data_out_349,
	output [15:0] data_out_350,
	output [15:0] data_out_351,
	output [15:0] data_out_352,
	output [15:0] data_out_353,
	output [15:0] data_out_354,
	output [15:0] data_out_355,
	output [15:0] data_out_356,
	output [15:0] data_out_357,
	output [15:0] data_out_358,
	output [15:0] data_out_359,
	output [15:0] data_out_360,
	output [15:0] data_out_361,
	output [15:0] data_out_362,
	output [15:0] data_out_363,
	output [15:0] data_out_364,
	output [15:0] data_out_365,
	output [15:0] data_out_366,
	output [15:0] data_out_367,
	output [15:0] data_out_368,
	output [15:0] data_out_369,
	output [15:0] data_out_370,
	output [15:0] data_out_371,
	output [15:0] data_out_372,
	output [15:0] data_out_373,
	output [15:0] data_out_374,
	output [15:0] data_out_375,
	output [15:0] data_out_376,
	output [15:0] data_out_377,
	output [15:0] data_out_378,
	output [15:0] data_out_379,
	output [15:0] data_out_380,
	output [15:0] data_out_381,
	output [15:0] data_out_382,
	output [15:0] data_out_383,
	output [15:0] data_out_384,
	output [15:0] data_out_385,
	output [15:0] data_out_386,
	output [15:0] data_out_387,
	output [15:0] data_out_388,
	output [15:0] data_out_389,
	output [15:0] data_out_390,
	output [15:0] data_out_391,
	output [15:0] data_out_392,
	output [15:0] data_out_393,
	output [15:0] data_out_394,
	output [15:0] data_out_395,
	output [15:0] data_out_396,
	output [15:0] data_out_397,
	output [15:0] data_out_398,
	output [15:0] data_out_399,
	output [15:0] data_out_400,
	output [15:0] data_out_401,
	output [15:0] data_out_402,
	output [15:0] data_out_403,
	output [15:0] data_out_404,
	output [15:0] data_out_405,
	output [15:0] data_out_406,
	output [15:0] data_out_407,
	output [15:0] data_out_408,
	output [15:0] data_out_409,
	output [15:0] data_out_410,
	output [15:0] data_out_411,
	output [15:0] data_out_412,
	output [15:0] data_out_413,
	output [15:0] data_out_414,
	output [15:0] data_out_415,
	output [15:0] data_out_416,
	output [15:0] data_out_417,
	output [15:0] data_out_418,
	output [15:0] data_out_419,
	output [15:0] data_out_420,
	output [15:0] data_out_421,
	output [15:0] data_out_422,
	output [15:0] data_out_423,
	output [15:0] data_out_424,
	output [15:0] data_out_425,
	output [15:0] data_out_426,
	output [15:0] data_out_427,
	output [15:0] data_out_428,
	output [15:0] data_out_429,
	output [15:0] data_out_430,
	output [15:0] data_out_431,
	output [15:0] data_out_432,
	output [15:0] data_out_433,
	output [15:0] data_out_434,
	output [15:0] data_out_435,
	output [15:0] data_out_436,
	output [15:0] data_out_437,
	output [15:0] data_out_438,
	output [15:0] data_out_439,
	output [15:0] data_out_440,
	output [15:0] data_out_441,
	output [15:0] data_out_442,
	output [15:0] data_out_443,
	output [15:0] data_out_444,
	output [15:0] data_out_445,
	output [15:0] data_out_446,
	output [15:0] data_out_447,
	output [15:0] data_out_448,
	output [15:0] data_out_449,
	output [15:0] data_out_450,
	output [15:0] data_out_451,
	output [15:0] data_out_452,
	output [15:0] data_out_453,
	output [15:0] data_out_454,
	output [15:0] data_out_455,
	output [15:0] data_out_456,
	output [15:0] data_out_457,
	output [15:0] data_out_458,
	output [15:0] data_out_459,
	output [15:0] data_out_460,
	output [15:0] data_out_461,
	output [15:0] data_out_462,
	output [15:0] data_out_463,
	output [15:0] data_out_464,
	output [15:0] data_out_465,
	output [15:0] data_out_466,
	output [15:0] data_out_467,
	output [15:0] data_out_468,
	output [15:0] data_out_469,
	output [15:0] data_out_470,
	output [15:0] data_out_471,
	output [15:0] data_out_472,
	output [15:0] data_out_473,
	output [15:0] data_out_474,
	output [15:0] data_out_475,
	output [15:0] data_out_476,
	output [15:0] data_out_477,
	output [15:0] data_out_478,
	output [15:0] data_out_479,
	output [15:0] data_out_480,
	output [15:0] data_out_481,
	output [15:0] data_out_482,
	output [15:0] data_out_483,
	output [15:0] data_out_484,
	output [15:0] data_out_485,
	output [15:0] data_out_486,
	output [15:0] data_out_487,
	output [15:0] data_out_488,
	output [15:0] data_out_489,
	output [15:0] data_out_490,
	output [15:0] data_out_491,
	output [15:0] data_out_492,
	output [15:0] data_out_493,
	output [15:0] data_out_494,
	output [15:0] data_out_495,
	output [15:0] data_out_496,
	output [15:0] data_out_497,
	output [15:0] data_out_498,
	output [15:0] data_out_499,
	output [15:0] data_out_500,
	output [15:0] data_out_501,
	output [15:0] data_out_502,
	output [15:0] data_out_503,
	output [15:0] data_out_504,
	output [15:0] data_out_505,
	output [15:0] data_out_506,
	output [15:0] data_out_507,
	output [15:0] data_out_508,
	output [15:0] data_out_509,
	output [15:0] data_out_510,
	output [15:0] data_out_511,
	output [15:0] data_out_512,
	output [15:0] data_out_513,
	output [15:0] data_out_514,
	output [15:0] data_out_515,
	output [15:0] data_out_516,
	output [15:0] data_out_517,
	output [15:0] data_out_518,
	output [15:0] data_out_519,
	output [15:0] data_out_520,
	output [15:0] data_out_521,
	output [15:0] data_out_522,
	output [15:0] data_out_523,
	output [15:0] data_out_524,
	output [15:0] data_out_525,
	output [15:0] data_out_526,
	output [15:0] data_out_527,
	output [15:0] data_out_528,
	output [15:0] data_out_529,
	output [15:0] data_out_530,
	output [15:0] data_out_531,
	output [15:0] data_out_532,
	output [15:0] data_out_533,
	output [15:0] data_out_534,
	output [15:0] data_out_535,
	output [15:0] data_out_536,
	output [15:0] data_out_537,
	output [15:0] data_out_538,
	output [15:0] data_out_539,
	output [15:0] data_out_540,
	output [15:0] data_out_541,
	output [15:0] data_out_542,
	output [15:0] data_out_543,
	output [15:0] data_out_544,
	output [15:0] data_out_545,
	output [15:0] data_out_546,
	output [15:0] data_out_547,
	output [15:0] data_out_548,
	output [15:0] data_out_549,
	output [15:0] data_out_550,
	output [15:0] data_out_551,
	output [15:0] data_out_552,
	output [15:0] data_out_553,
	output [15:0] data_out_554,
	output [15:0] data_out_555,
	output [15:0] data_out_556,
	output [15:0] data_out_557,
	output [15:0] data_out_558,
	output [15:0] data_out_559,
	output [15:0] data_out_560,
	output [15:0] data_out_561,
	output [15:0] data_out_562,
	output [15:0] data_out_563,
	output [15:0] data_out_564,
	output [15:0] data_out_565,
	output [15:0] data_out_566,
	output [15:0] data_out_567,
	output [15:0] data_out_568,
	output [15:0] data_out_569,
	output [15:0] data_out_570,
	output [15:0] data_out_571,
	output [15:0] data_out_572,
	output [15:0] data_out_573,
	output [15:0] data_out_574,
	output [15:0] data_out_575,
	output [15:0] data_out_576,
	output [15:0] data_out_577,
	output [15:0] data_out_578,
	output [15:0] data_out_579,
	output [15:0] data_out_580,
	output [15:0] data_out_581,
	output [15:0] data_out_582,
	output [15:0] data_out_583,
	output [15:0] data_out_584,
	output [15:0] data_out_585,
	output [15:0] data_out_586,
	output [15:0] data_out_587,
	output [15:0] data_out_588,
	output [15:0] data_out_589,
	output [15:0] data_out_590,
	output [15:0] data_out_591,
	output [15:0] data_out_592,
	output [15:0] data_out_593,
	output [15:0] data_out_594,
	output [15:0] data_out_595,
	output [15:0] data_out_596,
	output [15:0] data_out_597,
	output [15:0] data_out_598,
	output [15:0] data_out_599,
	output [15:0] data_out_600,
	output [15:0] data_out_601,
	output [15:0] data_out_602,
	output [15:0] data_out_603,
	output [15:0] data_out_604,
	output [15:0] data_out_605,
	output [15:0] data_out_606,
	output [15:0] data_out_607,
	output [15:0] data_out_608,
	output [15:0] data_out_609,
	output [15:0] data_out_610,
	output [15:0] data_out_611,
	output [15:0] data_out_612,
	output [15:0] data_out_613,
	output [15:0] data_out_614,
	output [15:0] data_out_615,
	output [15:0] data_out_616,
	output [15:0] data_out_617,
	output [15:0] data_out_618,
	output [15:0] data_out_619,
	output [15:0] data_out_620,
	output [15:0] data_out_621,
	output [15:0] data_out_622,
	output [15:0] data_out_623,
	output [15:0] data_out_624,
	output [15:0] data_out_625,
	output [15:0] data_out_626,
	output [15:0] data_out_627,
	output [15:0] data_out_628,
	output [15:0] data_out_629,
	output [15:0] data_out_630,
	output [15:0] data_out_631,
	output [15:0] data_out_632,
	output [15:0] data_out_633,
	output [15:0] data_out_634,
	output [15:0] data_out_635,
	output [15:0] data_out_636,
	output [15:0] data_out_637,
	output [15:0] data_out_638,
	output [15:0] data_out_639,
	output [15:0] data_out_640,
	output [15:0] data_out_641,
	output [15:0] data_out_642,
	output [15:0] data_out_643,
	output [15:0] data_out_644,
	output [15:0] data_out_645,
	output [15:0] data_out_646,
	output [15:0] data_out_647,
	output [15:0] data_out_648,
	output [15:0] data_out_649,
	output [15:0] data_out_650,
	output [15:0] data_out_651,
	output [15:0] data_out_652,
	output [15:0] data_out_653,
	output [15:0] data_out_654,
	output [15:0] data_out_655,
	output [15:0] data_out_656,
	output [15:0] data_out_657,
	output [15:0] data_out_658,
	output [15:0] data_out_659,
	output [15:0] data_out_660,
	output [15:0] data_out_661,
	output [15:0] data_out_662,
	output [15:0] data_out_663,
	output [15:0] data_out_664,
	output [15:0] data_out_665,
	output [15:0] data_out_666,
	output [15:0] data_out_667,
	output [15:0] data_out_668,
	output [15:0] data_out_669,
	output [15:0] data_out_670,
	output [15:0] data_out_671,
	output [15:0] data_out_672,
	output [15:0] data_out_673,
	output [15:0] data_out_674,
	output [15:0] data_out_675,
	output [15:0] data_out_676,
	output [15:0] data_out_677,
	output [15:0] data_out_678,
	output [15:0] data_out_679,
	output [15:0] data_out_680,
	output [15:0] data_out_681,
	output [15:0] data_out_682,
	output [15:0] data_out_683,
	output [15:0] data_out_684,
	output [15:0] data_out_685,
	output [15:0] data_out_686,
	output [15:0] data_out_687,
	output [15:0] data_out_688,
	output [15:0] data_out_689,
	output [15:0] data_out_690,
	output [15:0] data_out_691,
	output [15:0] data_out_692,
	output [15:0] data_out_693,
	output [15:0] data_out_694,
	output [15:0] data_out_695,
	output [15:0] data_out_696,
	output [15:0] data_out_697,
	output [15:0] data_out_698,
	output [15:0] data_out_699,
	output [15:0] data_out_700,
	output [15:0] data_out_701,
	output [15:0] data_out_702,
	output [15:0] data_out_703,
	output [15:0] data_out_704,
	output [15:0] data_out_705,
	output [15:0] data_out_706,
	output [15:0] data_out_707,
	output [15:0] data_out_708,
	output [15:0] data_out_709,
	output [15:0] data_out_710,
	output [15:0] data_out_711,
	output [15:0] data_out_712,
	output [15:0] data_out_713,
	output [15:0] data_out_714,
	output [15:0] data_out_715,
	output [15:0] data_out_716,
	output [15:0] data_out_717,
	output [15:0] data_out_718,
	output [15:0] data_out_719,
	output [15:0] data_out_720,
	output [15:0] data_out_721,
	output [15:0] data_out_722,
	output [15:0] data_out_723,
	output [15:0] data_out_724,
	output [15:0] data_out_725,
	output [15:0] data_out_726,
	output [15:0] data_out_727,
	output [15:0] data_out_728,
	output [15:0] data_out_729,
	output [15:0] data_out_730,
	output [15:0] data_out_731,
	output [15:0] data_out_732,
	output [15:0] data_out_733,
	output [15:0] data_out_734,
	output [15:0] data_out_735,
	output [15:0] data_out_736,
	output [15:0] data_out_737,
	output [15:0] data_out_738,
	output [15:0] data_out_739

	
	
	
	
);

    // ROM data initialization (example weights for simplicity)
    // Define a 192 x 16-bit memory array
    (* ram_style = "block" *) reg [15:0] rom_data [0:739]; 
	
	// Preload memory from a file during initialization
    initial begin
        $readmemh("weight_rom.hex", rom_data);     // Load the instruction memory from the hex file
    end
	
			assign data_out_0  = rom_data[0];
			assign data_out_1  = rom_data[1];
			assign data_out_2  = rom_data[2];
			assign data_out_3  = rom_data[3];
			assign data_out_4  = rom_data[4];
			assign data_out_5  = rom_data[5];
			assign data_out_6  = rom_data[6];
			assign data_out_7  = rom_data[7];
			assign data_out_8  = rom_data[8];
			assign data_out_9  = rom_data[9];
			assign data_out_10  = rom_data[10];
			assign data_out_11  = rom_data[11];
			assign data_out_12  = rom_data[12];
			assign data_out_13  = rom_data[13];
			assign data_out_14  = rom_data[14];
			assign data_out_15  = rom_data[15];
			assign data_out_16  = rom_data[16];
			assign data_out_17  = rom_data[17];
			assign data_out_18  = rom_data[18];
			assign data_out_19  = rom_data[19];
			assign data_out_20  = rom_data[20];
			assign data_out_21  = rom_data[21];
			assign data_out_22  = rom_data[22];
			assign data_out_23  = rom_data[23];
			assign data_out_24  = rom_data[24];
			assign data_out_25  = rom_data[25];
			assign data_out_26  = rom_data[26];
			assign data_out_27  = rom_data[27];
			assign data_out_28  = rom_data[28];
			assign data_out_29  = rom_data[29];
			assign data_out_30  = rom_data[30];
			assign data_out_31  = rom_data[31];
			assign data_out_32  = rom_data[32];
			assign data_out_33  = rom_data[33];
			assign data_out_34  = rom_data[34];
			assign data_out_35  = rom_data[35];
			assign data_out_36  = rom_data[36];
			assign data_out_37  = rom_data[37];
			assign data_out_38  = rom_data[38];
			assign data_out_39  = rom_data[39];
			assign data_out_40  = rom_data[40];
			assign data_out_41  = rom_data[41];
			assign data_out_42  = rom_data[42];
			assign data_out_43  = rom_data[43];
			assign data_out_44  = rom_data[44];
			assign data_out_45  = rom_data[45];
			assign data_out_46  = rom_data[46];
			assign data_out_47  = rom_data[47];
			assign data_out_48  = rom_data[48];
			assign data_out_49  = rom_data[49];
			assign data_out_50  = rom_data[50];
			assign data_out_51  = rom_data[51];
			assign data_out_52  = rom_data[52];
			assign data_out_53  = rom_data[53];
			assign data_out_54  = rom_data[54];
			assign data_out_55  = rom_data[55];
			assign data_out_56  = rom_data[56];
			assign data_out_57  = rom_data[57];
			assign data_out_58  = rom_data[58];
			assign data_out_59  = rom_data[59];
			assign data_out_60  = rom_data[60];
			assign data_out_61  = rom_data[61];
			assign data_out_62  = rom_data[62];
			assign data_out_63  = rom_data[63];
			assign data_out_64  = rom_data[64];
			assign data_out_65  = rom_data[65];
			assign data_out_66  = rom_data[66];
			assign data_out_67  = rom_data[67];
			assign data_out_68  = rom_data[68];
			assign data_out_69  = rom_data[69];
			assign data_out_70  = rom_data[70];
			assign data_out_71  = rom_data[71];
			assign data_out_72  = rom_data[72];
			assign data_out_73  = rom_data[73];
			assign data_out_74  = rom_data[74];
			assign data_out_75  = rom_data[75];
			assign data_out_76  = rom_data[76];
			assign data_out_77  = rom_data[77];
			assign data_out_78  = rom_data[78];
			assign data_out_79  = rom_data[79];
			assign data_out_80  = rom_data[80];
			assign data_out_81  = rom_data[81];
			assign data_out_82  = rom_data[82];
			assign data_out_83  = rom_data[83];
			assign data_out_84  = rom_data[84];
			assign data_out_85  = rom_data[85];
			assign data_out_86  = rom_data[86];
			assign data_out_87  = rom_data[87];
			assign data_out_88  = rom_data[88];
			assign data_out_89  = rom_data[89];
			assign data_out_90  = rom_data[90];
			assign data_out_91  = rom_data[91];
			assign data_out_92  = rom_data[92];
			assign data_out_93  = rom_data[93];
			assign data_out_94  = rom_data[94];
			assign data_out_95  = rom_data[95];
			assign data_out_96  = rom_data[96];
			assign data_out_97  = rom_data[97];
			assign data_out_98  = rom_data[98];
			assign data_out_99  = rom_data[99];
			assign data_out_100  = rom_data[100];
			assign data_out_101  = rom_data[101];
			assign data_out_102  = rom_data[102];
			assign data_out_103  = rom_data[103];
			assign data_out_104  = rom_data[104];
			assign data_out_105  = rom_data[105];
			assign data_out_106  = rom_data[106];
			assign data_out_107  = rom_data[107];
			assign data_out_108  = rom_data[108];
			assign data_out_109  = rom_data[109];
			assign data_out_110  = rom_data[110];
			assign data_out_111  = rom_data[111];
			assign data_out_112  = rom_data[112];
			assign data_out_113  = rom_data[113];
			assign data_out_114  = rom_data[114];
			assign data_out_115  = rom_data[115];
			assign data_out_116  = rom_data[116];
			assign data_out_117  = rom_data[117];
			assign data_out_118  = rom_data[118];
			assign data_out_119  = rom_data[119];
			assign data_out_120  = rom_data[120];
			assign data_out_121  = rom_data[121];
			assign data_out_122  = rom_data[122];
			assign data_out_123  = rom_data[123];
			assign data_out_124  = rom_data[124];
			assign data_out_125  = rom_data[125];
			assign data_out_126  = rom_data[126];
			assign data_out_127  = rom_data[127];
			assign data_out_128  = rom_data[128];
			assign data_out_129  = rom_data[129];
			assign data_out_130  = rom_data[130];
			assign data_out_131  = rom_data[131];
			assign data_out_132  = rom_data[132];
			assign data_out_133  = rom_data[133];
			assign data_out_134  = rom_data[134];
			assign data_out_135  = rom_data[135];
			assign data_out_136  = rom_data[136];
			assign data_out_137  = rom_data[137];
			assign data_out_138  = rom_data[138];
			assign data_out_139  = rom_data[139];
			assign data_out_140  = rom_data[140];
			assign data_out_141  = rom_data[141];
			assign data_out_142  = rom_data[142];
			assign data_out_143  = rom_data[143];
			assign data_out_144  = rom_data[144];
			assign data_out_145  = rom_data[145];
			assign data_out_146  = rom_data[146];
			assign data_out_147  = rom_data[147];
			assign data_out_148  = rom_data[148];
			assign data_out_149  = rom_data[149];
			assign data_out_150  = rom_data[150];
			assign data_out_151  = rom_data[151];
			assign data_out_152  = rom_data[152];
			assign data_out_153  = rom_data[153];
			assign data_out_154  = rom_data[154];
			assign data_out_155  = rom_data[155];
			assign data_out_156  = rom_data[156];
			assign data_out_157  = rom_data[157];
			assign data_out_158  = rom_data[158];
			assign data_out_159  = rom_data[159];
			assign data_out_160  = rom_data[160];
			assign data_out_161  = rom_data[161];
			assign data_out_162  = rom_data[162];
			assign data_out_163  = rom_data[163];
			assign data_out_164  = rom_data[164];
			assign data_out_165  = rom_data[165];
			assign data_out_166  = rom_data[166];
			assign data_out_167  = rom_data[167];
			assign data_out_168  = rom_data[168];
			assign data_out_169  = rom_data[169];
			assign data_out_170  = rom_data[170];
			assign data_out_171  = rom_data[171];
			assign data_out_172  = rom_data[172];
			assign data_out_173  = rom_data[173];
			assign data_out_174  = rom_data[174];
			assign data_out_175  = rom_data[175];
			assign data_out_176  = rom_data[176];
			assign data_out_177  = rom_data[177];
			assign data_out_178  = rom_data[178];
			assign data_out_179  = rom_data[179];
			assign data_out_180  = rom_data[180];
			assign data_out_181  = rom_data[181];
			assign data_out_182  = rom_data[182];
			assign data_out_183  = rom_data[183];
			assign data_out_184  = rom_data[184];
			assign data_out_185  = rom_data[185];
			assign data_out_186  = rom_data[186];
			assign data_out_187  = rom_data[187];
			assign data_out_188  = rom_data[188];
			assign data_out_189  = rom_data[189];
			assign data_out_190  = rom_data[190];
			assign data_out_191  = rom_data[191];
			assign data_out_192  = rom_data[192];
			assign data_out_193  = rom_data[193];
			assign data_out_194  = rom_data[194];
			assign data_out_195  = rom_data[195];
			assign data_out_196  = rom_data[196];
			assign data_out_197  = rom_data[197];
			assign data_out_198  = rom_data[198];
			assign data_out_199  = rom_data[199];
			assign data_out_200  = rom_data[200];
			assign data_out_201  = rom_data[201];
			assign data_out_202  = rom_data[202];
			assign data_out_203  = rom_data[203];
			assign data_out_204  = rom_data[204];
			assign data_out_205  = rom_data[205];
			assign data_out_206  = rom_data[206];
			assign data_out_207  = rom_data[207];
			assign data_out_208  = rom_data[208];
			assign data_out_209  = rom_data[209];
			assign data_out_210  = rom_data[210];
			assign data_out_211  = rom_data[211];
			assign data_out_212  = rom_data[212];
			assign data_out_213  = rom_data[213];
			assign data_out_214  = rom_data[214];
			assign data_out_215  = rom_data[215];
			assign data_out_216  = rom_data[216];
			assign data_out_217  = rom_data[217];
			assign data_out_218  = rom_data[218];
			assign data_out_219  = rom_data[219];
			assign data_out_220  = rom_data[220];
			assign data_out_221  = rom_data[221];
			assign data_out_222  = rom_data[222];
			assign data_out_223  = rom_data[223];
			assign data_out_224  = rom_data[224];
			assign data_out_225  = rom_data[225];
			assign data_out_226  = rom_data[226];
			assign data_out_227  = rom_data[227];
			assign data_out_228  = rom_data[228];
			assign data_out_229  = rom_data[229];
			assign data_out_230  = rom_data[230];
			assign data_out_231  = rom_data[231];
			assign data_out_232  = rom_data[232];
			assign data_out_233  = rom_data[233];
			assign data_out_234  = rom_data[234];
			assign data_out_235  = rom_data[235];
			assign data_out_236  = rom_data[236];
			assign data_out_237  = rom_data[237];
			assign data_out_238  = rom_data[238];
			assign data_out_239  = rom_data[239];
			assign data_out_240  = rom_data[240];
			assign data_out_241  = rom_data[241];
			assign data_out_242  = rom_data[242];
			assign data_out_243  = rom_data[243];
			assign data_out_244  = rom_data[244];
			assign data_out_245  = rom_data[245];
			assign data_out_246  = rom_data[246];
			assign data_out_247  = rom_data[247];
			assign data_out_248  = rom_data[248];
			assign data_out_249  = rom_data[249];
			assign data_out_250  = rom_data[250];
			assign data_out_251  = rom_data[251];
			assign data_out_252  = rom_data[252];
			assign data_out_253  = rom_data[253];
			assign data_out_254  = rom_data[254];
			assign data_out_255  = rom_data[255];
			assign data_out_256  = rom_data[256];
			assign data_out_257  = rom_data[257];
			assign data_out_258  = rom_data[258];
			assign data_out_259  = rom_data[259];
			assign data_out_260  = rom_data[260];
			assign data_out_261  = rom_data[261];
			assign data_out_262  = rom_data[262];
			assign data_out_263  = rom_data[263];
			assign data_out_264  = rom_data[264];
			assign data_out_265  = rom_data[265];
			assign data_out_266  = rom_data[266];
			assign data_out_267  = rom_data[267];
			assign data_out_268  = rom_data[268];
			assign data_out_269  = rom_data[269];
			assign data_out_270  = rom_data[270];
			assign data_out_271  = rom_data[271];
			assign data_out_272  = rom_data[272];
			assign data_out_273  = rom_data[273];
			assign data_out_274  = rom_data[274];
			assign data_out_275  = rom_data[275];
			assign data_out_276  = rom_data[276];
			assign data_out_277  = rom_data[277];
			assign data_out_278  = rom_data[278];
			assign data_out_279  = rom_data[279];
			assign data_out_280  = rom_data[280];
			assign data_out_281  = rom_data[281];
			assign data_out_282  = rom_data[282];
			assign data_out_283  = rom_data[283];
			assign data_out_284  = rom_data[284];
			assign data_out_285  = rom_data[285];
			assign data_out_286  = rom_data[286];
			assign data_out_287  = rom_data[287];
			assign data_out_288  = rom_data[288];
			assign data_out_289  = rom_data[289];
			assign data_out_290  = rom_data[290];
			assign data_out_291  = rom_data[291];
			assign data_out_292  = rom_data[292];
			assign data_out_293  = rom_data[293];
			assign data_out_294  = rom_data[294];
			assign data_out_295  = rom_data[295];
			assign data_out_296  = rom_data[296];
			assign data_out_297  = rom_data[297];
			assign data_out_298  = rom_data[298];
			assign data_out_299  = rom_data[299];
			assign data_out_300  = rom_data[300];
			assign data_out_301  = rom_data[301];
			assign data_out_302  = rom_data[302];
			assign data_out_303  = rom_data[303];
			assign data_out_304  = rom_data[304];
			assign data_out_305  = rom_data[305];
			assign data_out_306  = rom_data[306];
			assign data_out_307  = rom_data[307];
			assign data_out_308  = rom_data[308];
			assign data_out_309  = rom_data[309];
			assign data_out_310  = rom_data[310];
			assign data_out_311  = rom_data[311];
			assign data_out_312  = rom_data[312];
			assign data_out_313  = rom_data[313];
			assign data_out_314  = rom_data[314];
			assign data_out_315  = rom_data[315];
			assign data_out_316  = rom_data[316];
			assign data_out_317  = rom_data[317];
			assign data_out_318  = rom_data[318];
			assign data_out_319  = rom_data[319];
			assign data_out_320  = rom_data[320];
			assign data_out_321  = rom_data[321];
			assign data_out_322  = rom_data[322];
			assign data_out_323  = rom_data[323];
			assign data_out_324  = rom_data[324];
			assign data_out_325  = rom_data[325];
			assign data_out_326  = rom_data[326];
			assign data_out_327  = rom_data[327];
			assign data_out_328  = rom_data[328];
			assign data_out_329  = rom_data[329];
			assign data_out_330  = rom_data[330];
			assign data_out_331  = rom_data[331];
			assign data_out_332  = rom_data[332];
			assign data_out_333  = rom_data[333];
			assign data_out_334  = rom_data[334];
			assign data_out_335  = rom_data[335];
			assign data_out_336  = rom_data[336];
			assign data_out_337  = rom_data[337];
			assign data_out_338  = rom_data[338];
			assign data_out_339  = rom_data[339];
			assign data_out_340  = rom_data[340];
			assign data_out_341  = rom_data[341];
			assign data_out_342  = rom_data[342];
			assign data_out_343  = rom_data[343];
			assign data_out_344  = rom_data[344];
			assign data_out_345  = rom_data[345];
			assign data_out_346  = rom_data[346];
			assign data_out_347  = rom_data[347];
			assign data_out_348  = rom_data[348];
			assign data_out_349  = rom_data[349];
			assign data_out_350  = rom_data[350];
			assign data_out_351  = rom_data[351];
			assign data_out_352  = rom_data[352];
			assign data_out_353  = rom_data[353];
			assign data_out_354  = rom_data[354];
			assign data_out_355  = rom_data[355];
			assign data_out_356  = rom_data[356];
			assign data_out_357  = rom_data[357];
			assign data_out_358  = rom_data[358];
			assign data_out_359  = rom_data[359];
			assign data_out_360  = rom_data[360];
			assign data_out_361  = rom_data[361];
			assign data_out_362  = rom_data[362];
			assign data_out_363  = rom_data[363];
			assign data_out_364  = rom_data[364];
			assign data_out_365  = rom_data[365];
			assign data_out_366  = rom_data[366];
			assign data_out_367  = rom_data[367];
			assign data_out_368  = rom_data[368];
			assign data_out_369  = rom_data[369];
			assign data_out_370  = rom_data[370];
			assign data_out_371  = rom_data[371];
			assign data_out_372  = rom_data[372];
			assign data_out_373  = rom_data[373];
			assign data_out_374  = rom_data[374];
			assign data_out_375  = rom_data[375];
			assign data_out_376  = rom_data[376];
			assign data_out_377  = rom_data[377];
			assign data_out_378  = rom_data[378];
			assign data_out_379  = rom_data[379];
			assign data_out_380  = rom_data[380];
			assign data_out_381  = rom_data[381];
			assign data_out_382  = rom_data[382];
			assign data_out_383  = rom_data[383];
			assign data_out_384  = rom_data[384];
			assign data_out_385  = rom_data[385];
			assign data_out_386  = rom_data[386];
			assign data_out_387  = rom_data[387];
			assign data_out_388  = rom_data[388];
			assign data_out_389  = rom_data[389];
			assign data_out_390  = rom_data[390];
			assign data_out_391  = rom_data[391];
			assign data_out_392  = rom_data[392];
			assign data_out_393  = rom_data[393];
			assign data_out_394  = rom_data[394];
			assign data_out_395  = rom_data[395];
			assign data_out_396  = rom_data[396];
			assign data_out_397  = rom_data[397];
			assign data_out_398  = rom_data[398];
			assign data_out_399  = rom_data[399];
			assign data_out_400  = rom_data[400];
			assign data_out_401  = rom_data[401];
			assign data_out_402  = rom_data[402];
			assign data_out_403  = rom_data[403];
			assign data_out_404  = rom_data[404];
			assign data_out_405  = rom_data[405];
			assign data_out_406  = rom_data[406];
			assign data_out_407  = rom_data[407];
			assign data_out_408  = rom_data[408];
			assign data_out_409  = rom_data[409];
			assign data_out_410  = rom_data[410];
			assign data_out_411  = rom_data[411];
			assign data_out_412  = rom_data[412];
			assign data_out_413  = rom_data[413];
			assign data_out_414  = rom_data[414];
			assign data_out_415  = rom_data[415];
			assign data_out_416  = rom_data[416];
			assign data_out_417  = rom_data[417];
			assign data_out_418  = rom_data[418];
			assign data_out_419  = rom_data[419];
			assign data_out_420  = rom_data[420];
			assign data_out_421  = rom_data[421];
			assign data_out_422  = rom_data[422];
			assign data_out_423  = rom_data[423];
			assign data_out_424  = rom_data[424];
			assign data_out_425  = rom_data[425];
			assign data_out_426  = rom_data[426];
			assign data_out_427  = rom_data[427];
			assign data_out_428  = rom_data[428];
			assign data_out_429  = rom_data[429];
			assign data_out_430  = rom_data[430];
			assign data_out_431  = rom_data[431];
			assign data_out_432  = rom_data[432];
			assign data_out_433  = rom_data[433];
			assign data_out_434  = rom_data[434];
			assign data_out_435  = rom_data[435];
			assign data_out_436  = rom_data[436];
			assign data_out_437  = rom_data[437];
			assign data_out_438  = rom_data[438];
			assign data_out_439  = rom_data[439];
			assign data_out_440  = rom_data[440];
			assign data_out_441  = rom_data[441];
			assign data_out_442  = rom_data[442];
			assign data_out_443  = rom_data[443];
			assign data_out_444  = rom_data[444];
			assign data_out_445  = rom_data[445];
			assign data_out_446  = rom_data[446];
			assign data_out_447  = rom_data[447];
			assign data_out_448  = rom_data[448];
			assign data_out_449  = rom_data[449];
			assign data_out_450  = rom_data[450];
			assign data_out_451  = rom_data[451];
			assign data_out_452  = rom_data[452];
			assign data_out_453  = rom_data[453];
			assign data_out_454  = rom_data[454];
			assign data_out_455  = rom_data[455];
			assign data_out_456  = rom_data[456];
			assign data_out_457  = rom_data[457];
			assign data_out_458  = rom_data[458];
			assign data_out_459  = rom_data[459];
			assign data_out_460  = rom_data[460];
			assign data_out_461  = rom_data[461];
			assign data_out_462  = rom_data[462];
			assign data_out_463  = rom_data[463];
			assign data_out_464  = rom_data[464];
			assign data_out_465  = rom_data[465];
			assign data_out_466  = rom_data[466];
			assign data_out_467  = rom_data[467];
			assign data_out_468  = rom_data[468];
			assign data_out_469  = rom_data[469];
			assign data_out_470  = rom_data[470];
			assign data_out_471  = rom_data[471];
			assign data_out_472  = rom_data[472];
			assign data_out_473  = rom_data[473];
			assign data_out_474  = rom_data[474];
			assign data_out_475  = rom_data[475];
			assign data_out_476  = rom_data[476];
			assign data_out_477  = rom_data[477];
			assign data_out_478  = rom_data[478];
			assign data_out_479  = rom_data[479];
			assign data_out_480  = rom_data[480];
			assign data_out_481  = rom_data[481];
			assign data_out_482  = rom_data[482];
			assign data_out_483  = rom_data[483];
			assign data_out_484  = rom_data[484];
			assign data_out_485  = rom_data[485];
			assign data_out_486  = rom_data[486];
			assign data_out_487  = rom_data[487];
			assign data_out_488  = rom_data[488];
			assign data_out_489  = rom_data[489];
			assign data_out_490  = rom_data[490];
			assign data_out_491  = rom_data[491];
			assign data_out_492  = rom_data[492];
			assign data_out_493  = rom_data[493];
			assign data_out_494  = rom_data[494];
			assign data_out_495  = rom_data[495];
			assign data_out_496  = rom_data[496];
			assign data_out_497  = rom_data[497];
			assign data_out_498  = rom_data[498];
			assign data_out_499  = rom_data[499];
			assign data_out_500  = rom_data[500];
			assign data_out_501  = rom_data[501];
			assign data_out_502  = rom_data[502];
			assign data_out_503  = rom_data[503];
			assign data_out_504  = rom_data[504];
			assign data_out_505  = rom_data[505];
			assign data_out_506  = rom_data[506];
			assign data_out_507  = rom_data[507];
			assign data_out_508  = rom_data[508];
			assign data_out_509  = rom_data[509];
			assign data_out_510  = rom_data[510];
			assign data_out_511  = rom_data[511];
			assign data_out_512  = rom_data[512];
			assign data_out_513  = rom_data[513];
			assign data_out_514  = rom_data[514];
			assign data_out_515  = rom_data[515];
			assign data_out_516  = rom_data[516];
			assign data_out_517  = rom_data[517];
			assign data_out_518  = rom_data[518];
			assign data_out_519  = rom_data[519];
			assign data_out_520  = rom_data[520];
			assign data_out_521  = rom_data[521];
			assign data_out_522  = rom_data[522];
			assign data_out_523  = rom_data[523];
			assign data_out_524  = rom_data[524];
			assign data_out_525  = rom_data[525];
			assign data_out_526  = rom_data[526];
			assign data_out_527  = rom_data[527];
			assign data_out_528  = rom_data[528];
			assign data_out_529  = rom_data[529];
			assign data_out_530  = rom_data[530];
			assign data_out_531  = rom_data[531];
			assign data_out_532  = rom_data[532];
			assign data_out_533  = rom_data[533];
			assign data_out_534  = rom_data[534];
			assign data_out_535  = rom_data[535];
			assign data_out_536  = rom_data[536];
			assign data_out_537  = rom_data[537];
			assign data_out_538  = rom_data[538];
			assign data_out_539  = rom_data[539];
			assign data_out_540  = rom_data[540];
			assign data_out_541  = rom_data[541];
			assign data_out_542  = rom_data[542];
			assign data_out_543  = rom_data[543];
			assign data_out_544  = rom_data[544];
			assign data_out_545  = rom_data[545];
			assign data_out_546  = rom_data[546];
			assign data_out_547  = rom_data[547];
			assign data_out_548  = rom_data[548];
			assign data_out_549  = rom_data[549];
			assign data_out_550  = rom_data[550];
			assign data_out_551  = rom_data[551];
			assign data_out_552  = rom_data[552];
			assign data_out_553  = rom_data[553];
			assign data_out_554  = rom_data[554];
			assign data_out_555  = rom_data[555];
			assign data_out_556  = rom_data[556];
			assign data_out_557  = rom_data[557];
			assign data_out_558  = rom_data[558];
			assign data_out_559  = rom_data[559];
			assign data_out_560  = rom_data[560];
			assign data_out_561  = rom_data[561];
			assign data_out_562  = rom_data[562];
			assign data_out_563  = rom_data[563];
			assign data_out_564  = rom_data[564];
			assign data_out_565  = rom_data[565];
			assign data_out_566  = rom_data[566];
			assign data_out_567  = rom_data[567];
			assign data_out_568  = rom_data[568];
			assign data_out_569  = rom_data[569];
			assign data_out_570  = rom_data[570];
			assign data_out_571  = rom_data[571];
			assign data_out_572  = rom_data[572];
			assign data_out_573  = rom_data[573];
			assign data_out_574  = rom_data[574];
			assign data_out_575  = rom_data[575];
			assign data_out_576  = rom_data[576];
			assign data_out_577  = rom_data[577];
			assign data_out_578  = rom_data[578];
			assign data_out_579  = rom_data[579];
			assign data_out_580  = rom_data[580];
			assign data_out_581  = rom_data[581];
			assign data_out_582  = rom_data[582];
			assign data_out_583  = rom_data[583];
			assign data_out_584  = rom_data[584];
			assign data_out_585  = rom_data[585];
			assign data_out_586  = rom_data[586];
			assign data_out_587  = rom_data[587];
			assign data_out_588  = rom_data[588];
			assign data_out_589  = rom_data[589];
			assign data_out_590  = rom_data[590];
			assign data_out_591  = rom_data[591];
			assign data_out_592  = rom_data[592];
			assign data_out_593  = rom_data[593];
			assign data_out_594  = rom_data[594];
			assign data_out_595  = rom_data[595];
			assign data_out_596  = rom_data[596];
			assign data_out_597  = rom_data[597];
			assign data_out_598  = rom_data[598];
			assign data_out_599  = rom_data[599];
			assign data_out_600  = rom_data[600];
			assign data_out_601  = rom_data[601];
			assign data_out_602  = rom_data[602];
			assign data_out_603  = rom_data[603];
			assign data_out_604  = rom_data[604];
			assign data_out_605  = rom_data[605];
			assign data_out_606  = rom_data[606];
			assign data_out_607  = rom_data[607];
			assign data_out_608  = rom_data[608];
			assign data_out_609  = rom_data[609];
			assign data_out_610  = rom_data[610];
			assign data_out_611  = rom_data[611];
			assign data_out_612  = rom_data[612];
			assign data_out_613  = rom_data[613];
			assign data_out_614  = rom_data[614];
			assign data_out_615  = rom_data[615];
			assign data_out_616  = rom_data[616];
			assign data_out_617  = rom_data[617];
			assign data_out_618  = rom_data[618];
			assign data_out_619  = rom_data[619];
			assign data_out_620  = rom_data[620];
			assign data_out_621  = rom_data[621];
			assign data_out_622  = rom_data[622];
			assign data_out_623  = rom_data[623];
			assign data_out_624  = rom_data[624];
			assign data_out_625  = rom_data[625];
			assign data_out_626  = rom_data[626];
			assign data_out_627  = rom_data[627];
			assign data_out_628  = rom_data[628];
			assign data_out_629  = rom_data[629];
			assign data_out_630  = rom_data[630];
			assign data_out_631  = rom_data[631];
			assign data_out_632  = rom_data[632];
			assign data_out_633  = rom_data[633];
			assign data_out_634  = rom_data[634];
			assign data_out_635  = rom_data[635];
			assign data_out_636  = rom_data[636];
			assign data_out_637  = rom_data[637];
			assign data_out_638  = rom_data[638];
			assign data_out_639  = rom_data[639];
			assign data_out_640  = rom_data[640];
			assign data_out_641  = rom_data[641];
			assign data_out_642  = rom_data[642];
			assign data_out_643  = rom_data[643];
			assign data_out_644  = rom_data[644];
			assign data_out_645  = rom_data[645];
			assign data_out_646  = rom_data[646];
			assign data_out_647  = rom_data[647];
			assign data_out_648  = rom_data[648];
			assign data_out_649  = rom_data[649];
			assign data_out_650  = rom_data[650];
			assign data_out_651  = rom_data[651];
			assign data_out_652  = rom_data[652];
			assign data_out_653  = rom_data[653];
			assign data_out_654  = rom_data[654];
			assign data_out_655  = rom_data[655];
			assign data_out_656  = rom_data[656];
			assign data_out_657  = rom_data[657];
			assign data_out_658  = rom_data[658];
			assign data_out_659  = rom_data[659];
			assign data_out_660  = rom_data[660];
			assign data_out_661  = rom_data[661];
			assign data_out_662  = rom_data[662];
			assign data_out_663  = rom_data[663];
			assign data_out_664  = rom_data[664];
			assign data_out_665  = rom_data[665];
			assign data_out_666  = rom_data[666];
			assign data_out_667  = rom_data[667];
			assign data_out_668  = rom_data[668];
			assign data_out_669  = rom_data[669];
			assign data_out_670  = rom_data[670];
			assign data_out_671  = rom_data[671];
			assign data_out_672  = rom_data[672];
			assign data_out_673  = rom_data[673];
			assign data_out_674  = rom_data[674];
			assign data_out_675  = rom_data[675];
			assign data_out_676  = rom_data[676];
			assign data_out_677  = rom_data[677];
			assign data_out_678  = rom_data[678];
			assign data_out_679  = rom_data[679];
			assign data_out_680  = rom_data[680];
			assign data_out_681  = rom_data[681];
			assign data_out_682  = rom_data[682];
			assign data_out_683  = rom_data[683];
			assign data_out_684  = rom_data[684];
			assign data_out_685  = rom_data[685];
			assign data_out_686  = rom_data[686];
			assign data_out_687  = rom_data[687];
			assign data_out_688  = rom_data[688];
			assign data_out_689  = rom_data[689];
			assign data_out_690  = rom_data[690];
			assign data_out_691  = rom_data[691];
			assign data_out_692  = rom_data[692];
			assign data_out_693  = rom_data[693];
			assign data_out_694  = rom_data[694];
			assign data_out_695  = rom_data[695];
			assign data_out_696  = rom_data[696];
			assign data_out_697  = rom_data[697];
			assign data_out_698  = rom_data[698];
			assign data_out_699  = rom_data[699];
			assign data_out_700  = rom_data[700];
			assign data_out_701  = rom_data[701];
			assign data_out_702  = rom_data[702];
			assign data_out_703  = rom_data[703];
			assign data_out_704  = rom_data[704];
			assign data_out_705  = rom_data[705];
			assign data_out_706  = rom_data[706];
			assign data_out_707  = rom_data[707];
			assign data_out_708  = rom_data[708];
			assign data_out_709  = rom_data[709];
			assign data_out_710  = rom_data[710];
			assign data_out_711  = rom_data[711];
			assign data_out_712  = rom_data[712];
			assign data_out_713  = rom_data[713];
			assign data_out_714  = rom_data[714];
			assign data_out_715  = rom_data[715];
			assign data_out_716  = rom_data[716];
			assign data_out_717  = rom_data[717];
			assign data_out_718  = rom_data[718];
			assign data_out_719  = rom_data[719];
			assign data_out_720  = rom_data[720];
			assign data_out_721  = rom_data[721];
			assign data_out_722  = rom_data[722];
			assign data_out_723  = rom_data[723];
			assign data_out_724  = rom_data[724];
			assign data_out_725  = rom_data[725];
			assign data_out_726  = rom_data[726];
			assign data_out_727  = rom_data[727];
			assign data_out_728  = rom_data[728];
			assign data_out_729  = rom_data[729];
			assign data_out_730  = rom_data[730];
			assign data_out_731  = rom_data[731];
			assign data_out_732  = rom_data[732];
			assign data_out_733  = rom_data[733];
			assign data_out_734  = rom_data[734];
			assign data_out_735  = rom_data[735];
			assign data_out_736  = rom_data[736];
			assign data_out_737  = rom_data[737];
			assign data_out_738  = rom_data[738];
			assign data_out_739  = rom_data[739];


endmodule
