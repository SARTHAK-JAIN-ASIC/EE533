module weight_rom (
    input clk,
    input reset,
    output reg [15:0] data_out_0,
	output reg [15:0] data_out_1,
	output reg [15:0] data_out_2,
	output reg [15:0] data_out_3,
	output reg [15:0] data_out_4,
	output reg [15:0] data_out_5,
	output reg [15:0] data_out_6,
	output reg [15:0] data_out_7,
	output reg [15:0] data_out_8,
	output reg [15:0] data_out_9,
	output reg [15:0] data_out_10,
	output reg [15:0] data_out_11,
	output reg [15:0] data_out_12,
	output reg [15:0] data_out_13,
	output reg [15:0] data_out_14,
	output reg [15:0] data_out_15,
	output reg [15:0] data_out_16,
	output reg [15:0] data_out_17,
	output reg [15:0] data_out_18,
	output reg [15:0] data_out_19,
	output reg [15:0] data_out_20,
	output reg [15:0] data_out_21,
	output reg [15:0] data_out_22,
	output reg [15:0] data_out_23,
	output reg [15:0] data_out_24,
	output reg [15:0] data_out_25,
	output reg [15:0] data_out_26,
	output reg [15:0] data_out_27,
	output reg [15:0] data_out_28,
	output reg [15:0] data_out_29,
	output reg [15:0] data_out_30,
	output reg [15:0] data_out_31,
	output reg [15:0] data_out_32,
	output reg [15:0] data_out_33,
	output reg [15:0] data_out_34,
	output reg [15:0] data_out_35,
	output reg [15:0] data_out_36,
	output reg [15:0] data_out_37,
	output reg [15:0] data_out_38,
	output reg [15:0] data_out_39,
	output reg [15:0] data_out_40,
	output reg [15:0] data_out_41,
	output reg [15:0] data_out_42,
	output reg [15:0] data_out_43,
	output reg [15:0] data_out_44,
	output reg [15:0] data_out_45,
	output reg [15:0] data_out_46,
	output reg [15:0] data_out_47,
	output reg [15:0] data_out_48,
	output reg [15:0] data_out_49,
	output reg [15:0] data_out_50,
	output reg [15:0] data_out_51,
	output reg [15:0] data_out_52,
	output reg [15:0] data_out_53,
	output reg [15:0] data_out_54,
	output reg [15:0] data_out_55,
	output reg [15:0] data_out_56,
	output reg [15:0] data_out_57,
	output reg [15:0] data_out_58,
	output reg [15:0] data_out_59,
	output reg [15:0] data_out_60,
	output reg [15:0] data_out_61,
	output reg [15:0] data_out_62,
	output reg [15:0] data_out_63,
	output reg [15:0] data_out_64,
	output reg [15:0] data_out_65,
	output reg [15:0] data_out_66,
	output reg [15:0] data_out_67,
	output reg [15:0] data_out_68,
	output reg [15:0] data_out_69,
	output reg [15:0] data_out_70,
	output reg [15:0] data_out_71,
	output reg [15:0] data_out_72,
	output reg [15:0] data_out_73,
	output reg [15:0] data_out_74,
	output reg [15:0] data_out_75,
	output reg [15:0] data_out_76,
	output reg [15:0] data_out_77,
	output reg [15:0] data_out_78,
	output reg [15:0] data_out_79,
	output reg [15:0] data_out_80,
	output reg [15:0] data_out_81,
	output reg [15:0] data_out_82,
	output reg [15:0] data_out_83,
	output reg [15:0] data_out_84,
	output reg [15:0] data_out_85,
	output reg [15:0] data_out_86,
	output reg [15:0] data_out_87,
	output reg [15:0] data_out_88,
	output reg [15:0] data_out_89,
	output reg [15:0] data_out_90,
	output reg [15:0] data_out_91,
	output reg [15:0] data_out_92,
	output reg [15:0] data_out_93,
	output reg [15:0] data_out_94,
	output reg [15:0] data_out_95,
	output reg [15:0] data_out_96,
	output reg [15:0] data_out_97,
	output reg [15:0] data_out_98,
	output reg [15:0] data_out_99,
	output reg [15:0] data_out_100,
	output reg [15:0] data_out_101,
	output reg [15:0] data_out_102,
	output reg [15:0] data_out_103,
	output reg [15:0] data_out_104,
	output reg [15:0] data_out_105,
	output reg [15:0] data_out_106,
	output reg [15:0] data_out_107,
	output reg [15:0] data_out_108,
	output reg [15:0] data_out_109,
	output reg [15:0] data_out_110,
	output reg [15:0] data_out_111,
	output reg [15:0] data_out_112,
	output reg [15:0] data_out_113,
	output reg [15:0] data_out_114,
	output reg [15:0] data_out_115,
	output reg [15:0] data_out_116,
	output reg [15:0] data_out_117,
	output reg [15:0] data_out_118,
	output reg [15:0] data_out_119,
	output reg [15:0] data_out_120,
	output reg [15:0] data_out_121,
	output reg [15:0] data_out_122,
	output reg [15:0] data_out_123,
	output reg [15:0] data_out_124,
	output reg [15:0] data_out_125,
	output reg [15:0] data_out_126,
	output reg [15:0] data_out_127,
	output reg [15:0] data_out_128,
	output reg [15:0] data_out_129,
	output reg [15:0] data_out_130,
	output reg [15:0] data_out_131,
	output reg [15:0] data_out_132,
	output reg [15:0] data_out_133,
	output reg [15:0] data_out_134,
	output reg [15:0] data_out_135,
	output reg [15:0] data_out_136,
	output reg [15:0] data_out_137,
	output reg [15:0] data_out_138,
	output reg [15:0] data_out_139,
	output reg [15:0] data_out_140,
	output reg [15:0] data_out_141,
	output reg [15:0] data_out_142,
	output reg [15:0] data_out_143,
	output reg [15:0] data_out_144,
	output reg [15:0] data_out_145,
	output reg [15:0] data_out_146,
	output reg [15:0] data_out_147,
	output reg [15:0] data_out_148,
	output reg [15:0] data_out_149,
	output reg [15:0] data_out_150,
	output reg [15:0] data_out_151,
	output reg [15:0] data_out_152,
	output reg [15:0] data_out_153,
	output reg [15:0] data_out_154,
	output reg [15:0] data_out_155,
	output reg [15:0] data_out_156,
	output reg [15:0] data_out_157,
	output reg [15:0] data_out_158,
	output reg [15:0] data_out_159,
	output reg [15:0] data_out_160,
	output reg [15:0] data_out_161,
	output reg [15:0] data_out_162,
	output reg [15:0] data_out_163,
	output reg [15:0] data_out_164,
	output reg [15:0] data_out_165,
	output reg [15:0] data_out_166,
	output reg [15:0] data_out_167,
	output reg [15:0] data_out_168,
	output reg [15:0] data_out_169,
	output reg [15:0] data_out_170,
	output reg [15:0] data_out_171,
	output reg [15:0] data_out_172,
	output reg [15:0] data_out_173,
	output reg [15:0] data_out_174,
	output reg [15:0] data_out_175,
	output reg [15:0] data_out_176,
	output reg [15:0] data_out_177,
	output reg [15:0] data_out_178,
	output reg [15:0] data_out_179,
	output reg [15:0] data_out_180,
	output reg [15:0] data_out_181,
	output reg [15:0] data_out_182,
	output reg [15:0] data_out_183,
	output reg [15:0] data_out_184,
	output reg [15:0] data_out_185,
	output reg [15:0] data_out_186,
	output reg [15:0] data_out_187,
	output reg [15:0] data_out_188,
	output reg [15:0] data_out_189,
	output reg [15:0] data_out_190,
	output reg [15:0] data_out_191,
	output reg [15:0] data_out_192,
	output reg [15:0] data_out_193,
	output reg [15:0] data_out_194,
	output reg [15:0] data_out_195,
	output reg [15:0] data_out_196,
	output reg [15:0] data_out_197,
	output reg [15:0] data_out_198,
	output reg [15:0] data_out_199,
	output reg [15:0] data_out_200,
	output reg [15:0] data_out_201,
	output reg [15:0] data_out_202,
	output reg [15:0] data_out_203,
	output reg [15:0] data_out_204,
	output reg [15:0] data_out_205,
	output reg [15:0] data_out_206,
	output reg [15:0] data_out_207,
	output reg [15:0] data_out_208,
	output reg [15:0] data_out_209,
	output reg [15:0] data_out_210,
	output reg [15:0] data_out_211,
	output reg [15:0] data_out_212,
	output reg [15:0] data_out_213,
	output reg [15:0] data_out_214,
	output reg [15:0] data_out_215,
	output reg [15:0] data_out_216,
	output reg [15:0] data_out_217,
	output reg [15:0] data_out_218,
	output reg [15:0] data_out_219,
	output reg [15:0] data_out_220,
	output reg [15:0] data_out_221,
	output reg [15:0] data_out_222,
	output reg [15:0] data_out_223,
	output reg [15:0] data_out_224,
	output reg [15:0] data_out_225,
	output reg [15:0] data_out_226,
	output reg [15:0] data_out_227,
	output reg [15:0] data_out_228,
	output reg [15:0] data_out_229,
	output reg [15:0] data_out_230,
	output reg [15:0] data_out_231,
	output reg [15:0] data_out_232,
	output reg [15:0] data_out_233,
	output reg [15:0] data_out_234,
	output reg [15:0] data_out_235,
	output reg [15:0] data_out_236,
	output reg [15:0] data_out_237,
	output reg [15:0] data_out_238,
	output reg [15:0] data_out_239,
	output reg [15:0] data_out_240,
	output reg [15:0] data_out_241,
	output reg [15:0] data_out_242,
	output reg [15:0] data_out_243,
	output reg [15:0] data_out_244,
	output reg [15:0] data_out_245,
	output reg [15:0] data_out_246,
	output reg [15:0] data_out_247,
	output reg [15:0] data_out_248,
	output reg [15:0] data_out_249,
	output reg [15:0] data_out_250,
	output reg [15:0] data_out_251,
	output reg [15:0] data_out_252,
	output reg [15:0] data_out_253,
	output reg [15:0] data_out_254,
	output reg [15:0] data_out_255,
	output reg [15:0] data_out_256,
	output reg [15:0] data_out_257,
	output reg [15:0] data_out_258,
	output reg [15:0] data_out_259,
	output reg [15:0] data_out_260,
	output reg [15:0] data_out_261,
	output reg [15:0] data_out_262,
	output reg [15:0] data_out_263,
	output reg [15:0] data_out_264,
	output reg [15:0] data_out_265,
	output reg [15:0] data_out_266,
	output reg [15:0] data_out_267,
	output reg [15:0] data_out_268,
	output reg [15:0] data_out_269,
	output reg [15:0] data_out_270,
	output reg [15:0] data_out_271,
	output reg [15:0] data_out_272,
	output reg [15:0] data_out_273,
	output reg [15:0] data_out_274,
	output reg [15:0] data_out_275,
	output reg [15:0] data_out_276,
	output reg [15:0] data_out_277,
	output reg [15:0] data_out_278,
	output reg [15:0] data_out_279,
	output reg [15:0] data_out_280,
	output reg [15:0] data_out_281,
	output reg [15:0] data_out_282,
	output reg [15:0] data_out_283,
	output reg [15:0] data_out_284,
	output reg [15:0] data_out_285,
	output reg [15:0] data_out_286,
	output reg [15:0] data_out_287,
	output reg [15:0] data_out_288,
	output reg [15:0] data_out_289,
	output reg [15:0] data_out_290,
	output reg [15:0] data_out_291,
	output reg [15:0] data_out_292,
	output reg [15:0] data_out_293,
	output reg [15:0] data_out_294,
	output reg [15:0] data_out_295,
	output reg [15:0] data_out_296,
	output reg [15:0] data_out_297,
	output reg [15:0] data_out_298,
	output reg [15:0] data_out_299,
	output reg [15:0] data_out_300,
	output reg [15:0] data_out_301,
	output reg [15:0] data_out_302,
	output reg [15:0] data_out_303,
	output reg [15:0] data_out_304,
	output reg [15:0] data_out_305,
	output reg [15:0] data_out_306,
	output reg [15:0] data_out_307,
	output reg [15:0] data_out_308,
	output reg [15:0] data_out_309,
	output reg [15:0] data_out_310,
	output reg [15:0] data_out_311,
	output reg [15:0] data_out_312,
	output reg [15:0] data_out_313,
	output reg [15:0] data_out_314,
	output reg [15:0] data_out_315,
	output reg [15:0] data_out_316,
	output reg [15:0] data_out_317,
	output reg [15:0] data_out_318,
	output reg [15:0] data_out_319,
	output reg [15:0] data_out_320,
	output reg [15:0] data_out_321,
	output reg [15:0] data_out_322,
	output reg [15:0] data_out_323,
	output reg [15:0] data_out_324,
	output reg [15:0] data_out_325,
	output reg [15:0] data_out_326,
	output reg [15:0] data_out_327,
	output reg [15:0] data_out_328,
	output reg [15:0] data_out_329,
	output reg [15:0] data_out_330,
	output reg [15:0] data_out_331,
	output reg [15:0] data_out_332,
	output reg [15:0] data_out_333,
	output reg [15:0] data_out_334,
	output reg [15:0] data_out_335,
	output reg [15:0] data_out_336,
	output reg [15:0] data_out_337,
	output reg [15:0] data_out_338,
	output reg [15:0] data_out_339,
	output reg [15:0] data_out_340,
	output reg [15:0] data_out_341,
	output reg [15:0] data_out_342,
	output reg [15:0] data_out_343,
	output reg [15:0] data_out_344,
	output reg [15:0] data_out_345,
	output reg [15:0] data_out_346,
	output reg [15:0] data_out_347,
	output reg [15:0] data_out_348,
	output reg [15:0] data_out_349,
	output reg [15:0] data_out_350,
	output reg [15:0] data_out_351,
	output reg [15:0] data_out_352,
	output reg [15:0] data_out_353,
	output reg [15:0] data_out_354,
	output reg [15:0] data_out_355,
	output reg [15:0] data_out_356,
	output reg [15:0] data_out_357,
	output reg [15:0] data_out_358,
	output reg [15:0] data_out_359,
	output reg [15:0] data_out_360,
	output reg [15:0] data_out_361,
	output reg [15:0] data_out_362,
	output reg [15:0] data_out_363,
	output reg [15:0] data_out_364,
	output reg [15:0] data_out_365,
	output reg [15:0] data_out_366,
	output reg [15:0] data_out_367,
	output reg [15:0] data_out_368,
	output reg [15:0] data_out_369,
	output reg [15:0] data_out_370,
	output reg [15:0] data_out_371,
	output reg [15:0] data_out_372,
	output reg [15:0] data_out_373,
	output reg [15:0] data_out_374,
	output reg [15:0] data_out_375,
	output reg [15:0] data_out_376,
	output reg [15:0] data_out_377,
	output reg [15:0] data_out_378,
	output reg [15:0] data_out_379,
	output reg [15:0] data_out_380,
	output reg [15:0] data_out_381,
	output reg [15:0] data_out_382,
	output reg [15:0] data_out_383,
	output reg [15:0] data_out_384,
	output reg [15:0] data_out_385,
	output reg [15:0] data_out_386,
	output reg [15:0] data_out_387,
	output reg [15:0] data_out_388,
	output reg [15:0] data_out_389,
	output reg [15:0] data_out_390,
	output reg [15:0] data_out_391,
	output reg [15:0] data_out_392,
	output reg [15:0] data_out_393,
	output reg [15:0] data_out_394,
	output reg [15:0] data_out_395,
	output reg [15:0] data_out_396,
	output reg [15:0] data_out_397,
	output reg [15:0] data_out_398,
	output reg [15:0] data_out_399,
	output reg [15:0] data_out_400,
	output reg [15:0] data_out_401,
	output reg [15:0] data_out_402,
	output reg [15:0] data_out_403,
	output reg [15:0] data_out_404,
	output reg [15:0] data_out_405,
	output reg [15:0] data_out_406,
	output reg [15:0] data_out_407,
	output reg [15:0] data_out_408,
	output reg [15:0] data_out_409,
	output reg [15:0] data_out_410,
	output reg [15:0] data_out_411,
	output reg [15:0] data_out_412,
	output reg [15:0] data_out_413,
	output reg [15:0] data_out_414,
	output reg [15:0] data_out_415,
	output reg [15:0] data_out_416,
	output reg [15:0] data_out_417,
	output reg [15:0] data_out_418,
	output reg [15:0] data_out_419,
	output reg [15:0] data_out_420,
	output reg [15:0] data_out_421,
	output reg [15:0] data_out_422,
	output reg [15:0] data_out_423,
	output reg [15:0] data_out_424,
	output reg [15:0] data_out_425,
	output reg [15:0] data_out_426,
	output reg [15:0] data_out_427,
	output reg [15:0] data_out_428,
	output reg [15:0] data_out_429,
	output reg [15:0] data_out_430,
	output reg [15:0] data_out_431,
	output reg [15:0] data_out_432,
	output reg [15:0] data_out_433,
	output reg [15:0] data_out_434,
	output reg [15:0] data_out_435,
	output reg [15:0] data_out_436,
	output reg [15:0] data_out_437,
	output reg [15:0] data_out_438,
	output reg [15:0] data_out_439,
	output reg [15:0] data_out_440,
	output reg [15:0] data_out_441,
	output reg [15:0] data_out_442,
	output reg [15:0] data_out_443,
	output reg [15:0] data_out_444,
	output reg [15:0] data_out_445,
	output reg [15:0] data_out_446,
	output reg [15:0] data_out_447,
	output reg [15:0] data_out_448,
	output reg [15:0] data_out_449,
	output reg [15:0] data_out_450,
	output reg [15:0] data_out_451,
	output reg [15:0] data_out_452,
	output reg [15:0] data_out_453,
	output reg [15:0] data_out_454,
	output reg [15:0] data_out_455,
	output reg [15:0] data_out_456,
	output reg [15:0] data_out_457,
	output reg [15:0] data_out_458,
	output reg [15:0] data_out_459,
	output reg [15:0] data_out_460,
	output reg [15:0] data_out_461,
	output reg [15:0] data_out_462,
	output reg [15:0] data_out_463,
	output reg [15:0] data_out_464,
	output reg [15:0] data_out_465,
	output reg [15:0] data_out_466,
	output reg [15:0] data_out_467,
	output reg [15:0] data_out_468,
	output reg [15:0] data_out_469,
	output reg [15:0] data_out_470,
	output reg [15:0] data_out_471,
	output reg [15:0] data_out_472,
	output reg [15:0] data_out_473,
	output reg [15:0] data_out_474,
	output reg [15:0] data_out_475,
	output reg [15:0] data_out_476,
	output reg [15:0] data_out_477,
	output reg [15:0] data_out_478,
	output reg [15:0] data_out_479,
	output reg [15:0] data_out_480,
	output reg [15:0] data_out_481,
	output reg [15:0] data_out_482,
	output reg [15:0] data_out_483,
	output reg [15:0] data_out_484,
	output reg [15:0] data_out_485,
	output reg [15:0] data_out_486,
	output reg [15:0] data_out_487,
	output reg [15:0] data_out_488,
	output reg [15:0] data_out_489,
	output reg [15:0] data_out_490,
	output reg [15:0] data_out_491,
	output reg [15:0] data_out_492,
	output reg [15:0] data_out_493,
	output reg [15:0] data_out_494,
	output reg [15:0] data_out_495,
	output reg [15:0] data_out_496,
	output reg [15:0] data_out_497,
	output reg [15:0] data_out_498,
	output reg [15:0] data_out_499,
	output reg [15:0] data_out_500,
	output reg [15:0] data_out_501,
	output reg [15:0] data_out_502,
	output reg [15:0] data_out_503,
	output reg [15:0] data_out_504,
	output reg [15:0] data_out_505,
	output reg [15:0] data_out_506,
	output reg [15:0] data_out_507,
	output reg [15:0] data_out_508,
	output reg [15:0] data_out_509,
	output reg [15:0] data_out_510,
	output reg [15:0] data_out_511,
	output reg [15:0] data_out_512,
	output reg [15:0] data_out_513,
	output reg [15:0] data_out_514,
	output reg [15:0] data_out_515,
	output reg [15:0] data_out_516,
	output reg [15:0] data_out_517,
	output reg [15:0] data_out_518,
	output reg [15:0] data_out_519,
	output reg [15:0] data_out_520,
	output reg [15:0] data_out_521,
	output reg [15:0] data_out_522,
	output reg [15:0] data_out_523,
	output reg [15:0] data_out_524,
	output reg [15:0] data_out_525,
	output reg [15:0] data_out_526,
	output reg [15:0] data_out_527,
	output reg [15:0] data_out_528,
	output reg [15:0] data_out_529,
	output reg [15:0] data_out_530,
	output reg [15:0] data_out_531,
	output reg [15:0] data_out_532,
	output reg [15:0] data_out_533,
	output reg [15:0] data_out_534,
	output reg [15:0] data_out_535,
	output reg [15:0] data_out_536,
	output reg [15:0] data_out_537,
	output reg [15:0] data_out_538,
	output reg [15:0] data_out_539,
	output reg [15:0] data_out_540,
	output reg [15:0] data_out_541,
	output reg [15:0] data_out_542,
	output reg [15:0] data_out_543,
	output reg [15:0] data_out_544,
	output reg [15:0] data_out_545,
	output reg [15:0] data_out_546,
	output reg [15:0] data_out_547,
	output reg [15:0] data_out_548,
	output reg [15:0] data_out_549,
	output reg [15:0] data_out_550,
	output reg [15:0] data_out_551,
	output reg [15:0] data_out_552,
	output reg [15:0] data_out_553,
	output reg [15:0] data_out_554,
	output reg [15:0] data_out_555,
	output reg [15:0] data_out_556,
	output reg [15:0] data_out_557,
	output reg [15:0] data_out_558,
	output reg [15:0] data_out_559,
	output reg [15:0] data_out_560,
	output reg [15:0] data_out_561,
	output reg [15:0] data_out_562,
	output reg [15:0] data_out_563,
	output reg [15:0] data_out_564,
	output reg [15:0] data_out_565,
	output reg [15:0] data_out_566,
	output reg [15:0] data_out_567,
	output reg [15:0] data_out_568,
	output reg [15:0] data_out_569,
	output reg [15:0] data_out_570,
	output reg [15:0] data_out_571,
	output reg [15:0] data_out_572,
	output reg [15:0] data_out_573,
	output reg [15:0] data_out_574,
	output reg [15:0] data_out_575,
	output reg [15:0] data_out_576,
	output reg [15:0] data_out_577,
	output reg [15:0] data_out_578,
	output reg [15:0] data_out_579,
	output reg [15:0] data_out_580,
	output reg [15:0] data_out_581,
	output reg [15:0] data_out_582,
	output reg [15:0] data_out_583,
	output reg [15:0] data_out_584,
	output reg [15:0] data_out_585,
	output reg [15:0] data_out_586,
	output reg [15:0] data_out_587,
	output reg [15:0] data_out_588,
	output reg [15:0] data_out_589,
	output reg [15:0] data_out_590,
	output reg [15:0] data_out_591,
	output reg [15:0] data_out_592,
	output reg [15:0] data_out_593,
	output reg [15:0] data_out_594,
	output reg [15:0] data_out_595,
	output reg [15:0] data_out_596,
	output reg [15:0] data_out_597,
	output reg [15:0] data_out_598,
	output reg [15:0] data_out_599,
	output reg [15:0] data_out_600,
	output reg [15:0] data_out_601,
	output reg [15:0] data_out_602,
	output reg [15:0] data_out_603,
	output reg [15:0] data_out_604,
	output reg [15:0] data_out_605,
	output reg [15:0] data_out_606,
	output reg [15:0] data_out_607,
	output reg [15:0] data_out_608,
	output reg [15:0] data_out_609,
	output reg [15:0] data_out_610,
	output reg [15:0] data_out_611,
	output reg [15:0] data_out_612,
	output reg [15:0] data_out_613,
	output reg [15:0] data_out_614,
	output reg [15:0] data_out_615,
	output reg [15:0] data_out_616,
	output reg [15:0] data_out_617,
	output reg [15:0] data_out_618,
	output reg [15:0] data_out_619,
	output reg [15:0] data_out_620,
	output reg [15:0] data_out_621,
	output reg [15:0] data_out_622,
	output reg [15:0] data_out_623,
	output reg [15:0] data_out_624,
	output reg [15:0] data_out_625,
	output reg [15:0] data_out_626,
	output reg [15:0] data_out_627,
	output reg [15:0] data_out_628,
	output reg [15:0] data_out_629,
	output reg [15:0] data_out_630,
	output reg [15:0] data_out_631,
	output reg [15:0] data_out_632,
	output reg [15:0] data_out_633,
	output reg [15:0] data_out_634,
	output reg [15:0] data_out_635,
	output reg [15:0] data_out_636,
	output reg [15:0] data_out_637,
	output reg [15:0] data_out_638,
	output reg [15:0] data_out_639,
	output reg [15:0] data_out_640,
	output reg [15:0] data_out_641,
	output reg [15:0] data_out_642,
	output reg [15:0] data_out_643,
	output reg [15:0] data_out_644,
	output reg [15:0] data_out_645,
	output reg [15:0] data_out_646,
	output reg [15:0] data_out_647,
	output reg [15:0] data_out_648,
	output reg [15:0] data_out_649,
	output reg [15:0] data_out_650,
	output reg [15:0] data_out_651,
	output reg [15:0] data_out_652,
	output reg [15:0] data_out_653,
	output reg [15:0] data_out_654,
	output reg [15:0] data_out_655,
	output reg [15:0] data_out_656,
	output reg [15:0] data_out_657,
	output reg [15:0] data_out_658,
	output reg [15:0] data_out_659,
	output reg [15:0] data_out_660,
	output reg [15:0] data_out_661,
	output reg [15:0] data_out_662,
	output reg [15:0] data_out_663,
	output reg [15:0] data_out_664,
	output reg [15:0] data_out_665,
	output reg [15:0] data_out_666,
	output reg [15:0] data_out_667,
	output reg [15:0] data_out_668,
	output reg [15:0] data_out_669,
	output reg [15:0] data_out_670,
	output reg [15:0] data_out_671,
	output reg [15:0] data_out_672,
	output reg [15:0] data_out_673,
	output reg [15:0] data_out_674,
	output reg [15:0] data_out_675,
	output reg [15:0] data_out_676,
	output reg [15:0] data_out_677,
	output reg [15:0] data_out_678,
	output reg [15:0] data_out_679,
	output reg [15:0] data_out_680,
	output reg [15:0] data_out_681,
	output reg [15:0] data_out_682,
	output reg [15:0] data_out_683,
	output reg [15:0] data_out_684,
	output reg [15:0] data_out_685,
	output reg [15:0] data_out_686,
	output reg [15:0] data_out_687,
	output reg [15:0] data_out_688,
	output reg [15:0] data_out_689,
	output reg [15:0] data_out_690,
	output reg [15:0] data_out_691,
	output reg [15:0] data_out_692,
	output reg [15:0] data_out_693,
	output reg [15:0] data_out_694,
	output reg [15:0] data_out_695,
	output reg [15:0] data_out_696,
	output reg [15:0] data_out_697,
	output reg [15:0] data_out_698,
	output reg [15:0] data_out_699,
	output reg [15:0] data_out_700,
	output reg [15:0] data_out_701,
	output reg [15:0] data_out_702,
	output reg [15:0] data_out_703,
	output reg [15:0] data_out_704,
	output reg [15:0] data_out_705,
	output reg [15:0] data_out_706,
	output reg [15:0] data_out_707,
	output reg [15:0] data_out_708,
	output reg [15:0] data_out_709,
	output reg [15:0] data_out_710,
	output reg [15:0] data_out_711,
	output reg [15:0] data_out_712,
	output reg [15:0] data_out_713,
	output reg [15:0] data_out_714,
	output reg [15:0] data_out_715,
	output reg [15:0] data_out_716,
	output reg [15:0] data_out_717,
	output reg [15:0] data_out_718,
	output reg [15:0] data_out_719,
	output reg [15:0] data_out_720,
	output reg [15:0] data_out_721,
	output reg [15:0] data_out_722,
	output reg [15:0] data_out_723,
	output reg [15:0] data_out_724,
	output reg [15:0] data_out_725,
	output reg [15:0] data_out_726,
	output reg [15:0] data_out_727,
	output reg [15:0] data_out_728,
	output reg [15:0] data_out_729,
	output reg [15:0] data_out_730,
	output reg [15:0] data_out_731,
	output reg [15:0] data_out_732,
	output reg [15:0] data_out_733,
	output reg [15:0] data_out_734,
	output reg [15:0] data_out_735,
	output reg [15:0] data_out_736,
	output reg [15:0] data_out_737,
	output reg [15:0] data_out_738,
	output reg [15:0] data_out_739

	
	
	
	
);

    // ROM data initialization (example weights for simplicity)
    // Define a 192 x 16-bit memory array
    (* ram_style = "block" *) reg [15:0] rom_data [0:739]; 
	
	// Preload memory from a file during initialization
    initial begin
        $readmemh("weight_rom.hex", rom_data);     // Load the instruction memory from the hex file
    end

    always @(posedge clk or posedge reset) begin
        if (reset) begin
            // Reset logic if needed
        end else begin
            // Fetch data from ROM based on the address
            data_out_0  <= rom_data[0];
			data_out_1  <= rom_data[1];
			data_out_2  <= rom_data[2];
			data_out_3  <= rom_data[3];
			data_out_4  <= rom_data[4];
			data_out_5  <= rom_data[5];
			data_out_6  <= rom_data[6];
			data_out_7  <= rom_data[7];
			data_out_8  <= rom_data[8];
			data_out_9  <= rom_data[9];
			data_out_10  <= rom_data[10];
			data_out_11  <= rom_data[11];
			data_out_12  <= rom_data[12];
			data_out_13  <= rom_data[13];
			data_out_14  <= rom_data[14];
			data_out_15  <= rom_data[15];
			data_out_16  <= rom_data[16];
			data_out_17  <= rom_data[17];
			data_out_18  <= rom_data[18];
			data_out_19  <= rom_data[19];
			data_out_20  <= rom_data[20];
			data_out_21  <= rom_data[21];
			data_out_22  <= rom_data[22];
			data_out_23  <= rom_data[23];
			data_out_24  <= rom_data[24];
			data_out_25  <= rom_data[25];
			data_out_26  <= rom_data[26];
			data_out_27  <= rom_data[27];
			data_out_28  <= rom_data[28];
			data_out_29  <= rom_data[29];
			data_out_30  <= rom_data[30];
			data_out_31  <= rom_data[31];
			data_out_32  <= rom_data[32];
			data_out_33  <= rom_data[33];
			data_out_34  <= rom_data[34];
			data_out_35  <= rom_data[35];
			data_out_36  <= rom_data[36];
			data_out_37  <= rom_data[37];
			data_out_38  <= rom_data[38];
			data_out_39  <= rom_data[39];
			data_out_40  <= rom_data[40];
			data_out_41  <= rom_data[41];
			data_out_42  <= rom_data[42];
			data_out_43  <= rom_data[43];
			data_out_44  <= rom_data[44];
			data_out_45  <= rom_data[45];
			data_out_46  <= rom_data[46];
			data_out_47  <= rom_data[47];
			data_out_48  <= rom_data[48];
			data_out_49  <= rom_data[49];
			data_out_50  <= rom_data[50];
			data_out_51  <= rom_data[51];
			data_out_52  <= rom_data[52];
			data_out_53  <= rom_data[53];
			data_out_54  <= rom_data[54];
			data_out_55  <= rom_data[55];
			data_out_56  <= rom_data[56];
			data_out_57  <= rom_data[57];
			data_out_58  <= rom_data[58];
			data_out_59  <= rom_data[59];
			data_out_60  <= rom_data[60];
			data_out_61  <= rom_data[61];
			data_out_62  <= rom_data[62];
			data_out_63  <= rom_data[63];
			data_out_64  <= rom_data[64];
			data_out_65  <= rom_data[65];
			data_out_66  <= rom_data[66];
			data_out_67  <= rom_data[67];
			data_out_68  <= rom_data[68];
			data_out_69  <= rom_data[69];
			data_out_70  <= rom_data[70];
			data_out_71  <= rom_data[71];
			data_out_72  <= rom_data[72];
			data_out_73  <= rom_data[73];
			data_out_74  <= rom_data[74];
			data_out_75  <= rom_data[75];
			data_out_76  <= rom_data[76];
			data_out_77  <= rom_data[77];
			data_out_78  <= rom_data[78];
			data_out_79  <= rom_data[79];
			data_out_80  <= rom_data[80];
			data_out_81  <= rom_data[81];
			data_out_82  <= rom_data[82];
			data_out_83  <= rom_data[83];
			data_out_84  <= rom_data[84];
			data_out_85  <= rom_data[85];
			data_out_86  <= rom_data[86];
			data_out_87  <= rom_data[87];
			data_out_88  <= rom_data[88];
			data_out_89  <= rom_data[89];
			data_out_90  <= rom_data[90];
			data_out_91  <= rom_data[91];
			data_out_92  <= rom_data[92];
			data_out_93  <= rom_data[93];
			data_out_94  <= rom_data[94];
			data_out_95  <= rom_data[95];
			data_out_96  <= rom_data[96];
			data_out_97  <= rom_data[97];
			data_out_98  <= rom_data[98];
			data_out_99  <= rom_data[99];
			data_out_100  <= rom_data[100];
			data_out_101  <= rom_data[101];
			data_out_102  <= rom_data[102];
			data_out_103  <= rom_data[103];
			data_out_104  <= rom_data[104];
			data_out_105  <= rom_data[105];
			data_out_106  <= rom_data[106];
			data_out_107  <= rom_data[107];
			data_out_108  <= rom_data[108];
			data_out_109  <= rom_data[109];
			data_out_110  <= rom_data[110];
			data_out_111  <= rom_data[111];
			data_out_112  <= rom_data[112];
			data_out_113  <= rom_data[113];
			data_out_114  <= rom_data[114];
			data_out_115  <= rom_data[115];
			data_out_116  <= rom_data[116];
			data_out_117  <= rom_data[117];
			data_out_118  <= rom_data[118];
			data_out_119  <= rom_data[119];
			data_out_120  <= rom_data[120];
			data_out_121  <= rom_data[121];
			data_out_122  <= rom_data[122];
			data_out_123  <= rom_data[123];
			data_out_124  <= rom_data[124];
			data_out_125  <= rom_data[125];
			data_out_126  <= rom_data[126];
			data_out_127  <= rom_data[127];
			data_out_128  <= rom_data[128];
			data_out_129  <= rom_data[129];
			data_out_130  <= rom_data[130];
			data_out_131  <= rom_data[131];
			data_out_132  <= rom_data[132];
			data_out_133  <= rom_data[133];
			data_out_134  <= rom_data[134];
			data_out_135  <= rom_data[135];
			data_out_136  <= rom_data[136];
			data_out_137  <= rom_data[137];
			data_out_138  <= rom_data[138];
			data_out_139  <= rom_data[139];
			data_out_140  <= rom_data[140];
			data_out_141  <= rom_data[141];
			data_out_142  <= rom_data[142];
			data_out_143  <= rom_data[143];
			data_out_144  <= rom_data[144];
			data_out_145  <= rom_data[145];
			data_out_146  <= rom_data[146];
			data_out_147  <= rom_data[147];
			data_out_148  <= rom_data[148];
			data_out_149  <= rom_data[149];
			data_out_150  <= rom_data[150];
			data_out_151  <= rom_data[151];
			data_out_152  <= rom_data[152];
			data_out_153  <= rom_data[153];
			data_out_154  <= rom_data[154];
			data_out_155  <= rom_data[155];
			data_out_156  <= rom_data[156];
			data_out_157  <= rom_data[157];
			data_out_158  <= rom_data[158];
			data_out_159  <= rom_data[159];
			data_out_160  <= rom_data[160];
			data_out_161  <= rom_data[161];
			data_out_162  <= rom_data[162];
			data_out_163  <= rom_data[163];
			data_out_164  <= rom_data[164];
			data_out_165  <= rom_data[165];
			data_out_166  <= rom_data[166];
			data_out_167  <= rom_data[167];
			data_out_168  <= rom_data[168];
			data_out_169  <= rom_data[169];
			data_out_170  <= rom_data[170];
			data_out_171  <= rom_data[171];
			data_out_172  <= rom_data[172];
			data_out_173  <= rom_data[173];
			data_out_174  <= rom_data[174];
			data_out_175  <= rom_data[175];
			data_out_176  <= rom_data[176];
			data_out_177  <= rom_data[177];
			data_out_178  <= rom_data[178];
			data_out_179  <= rom_data[179];
			data_out_180  <= rom_data[180];
			data_out_181  <= rom_data[181];
			data_out_182  <= rom_data[182];
			data_out_183  <= rom_data[183];
			data_out_184  <= rom_data[184];
			data_out_185  <= rom_data[185];
			data_out_186  <= rom_data[186];
			data_out_187  <= rom_data[187];
			data_out_188  <= rom_data[188];
			data_out_189  <= rom_data[189];
			data_out_190  <= rom_data[190];
			data_out_191  <= rom_data[191];
			data_out_192  <= rom_data[192];
			data_out_193  <= rom_data[193];
			data_out_194  <= rom_data[194];
			data_out_195  <= rom_data[195];
			data_out_196  <= rom_data[196];
			data_out_197  <= rom_data[197];
			data_out_198  <= rom_data[198];
			data_out_199  <= rom_data[199];
			data_out_200  <= rom_data[200];
			data_out_201  <= rom_data[201];
			data_out_202  <= rom_data[202];
			data_out_203  <= rom_data[203];
			data_out_204  <= rom_data[204];
			data_out_205  <= rom_data[205];
			data_out_206  <= rom_data[206];
			data_out_207  <= rom_data[207];
			data_out_208  <= rom_data[208];
			data_out_209  <= rom_data[209];
			data_out_210  <= rom_data[210];
			data_out_211  <= rom_data[211];
			data_out_212  <= rom_data[212];
			data_out_213  <= rom_data[213];
			data_out_214  <= rom_data[214];
			data_out_215  <= rom_data[215];
			data_out_216  <= rom_data[216];
			data_out_217  <= rom_data[217];
			data_out_218  <= rom_data[218];
			data_out_219  <= rom_data[219];
			data_out_220  <= rom_data[220];
			data_out_221  <= rom_data[221];
			data_out_222  <= rom_data[222];
			data_out_223  <= rom_data[223];
			data_out_224  <= rom_data[224];
			data_out_225  <= rom_data[225];
			data_out_226  <= rom_data[226];
			data_out_227  <= rom_data[227];
			data_out_228  <= rom_data[228];
			data_out_229  <= rom_data[229];
			data_out_230  <= rom_data[230];
			data_out_231  <= rom_data[231];
			data_out_232  <= rom_data[232];
			data_out_233  <= rom_data[233];
			data_out_234  <= rom_data[234];
			data_out_235  <= rom_data[235];
			data_out_236  <= rom_data[236];
			data_out_237  <= rom_data[237];
			data_out_238  <= rom_data[238];
			data_out_239  <= rom_data[239];
			data_out_240  <= rom_data[240];
			data_out_241  <= rom_data[241];
			data_out_242  <= rom_data[242];
			data_out_243  <= rom_data[243];
			data_out_244  <= rom_data[244];
			data_out_245  <= rom_data[245];
			data_out_246  <= rom_data[246];
			data_out_247  <= rom_data[247];
			data_out_248  <= rom_data[248];
			data_out_249  <= rom_data[249];
			data_out_250  <= rom_data[250];
			data_out_251  <= rom_data[251];
			data_out_252  <= rom_data[252];
			data_out_253  <= rom_data[253];
			data_out_254  <= rom_data[254];
			data_out_255  <= rom_data[255];
			data_out_256  <= rom_data[256];
			data_out_257  <= rom_data[257];
			data_out_258  <= rom_data[258];
			data_out_259  <= rom_data[259];
			data_out_260  <= rom_data[260];
			data_out_261  <= rom_data[261];
			data_out_262  <= rom_data[262];
			data_out_263  <= rom_data[263];
			data_out_264  <= rom_data[264];
			data_out_265  <= rom_data[265];
			data_out_266  <= rom_data[266];
			data_out_267  <= rom_data[267];
			data_out_268  <= rom_data[268];
			data_out_269  <= rom_data[269];
			data_out_270  <= rom_data[270];
			data_out_271  <= rom_data[271];
			data_out_272  <= rom_data[272];
			data_out_273  <= rom_data[273];
			data_out_274  <= rom_data[274];
			data_out_275  <= rom_data[275];
			data_out_276  <= rom_data[276];
			data_out_277  <= rom_data[277];
			data_out_278  <= rom_data[278];
			data_out_279  <= rom_data[279];
			data_out_280  <= rom_data[280];
			data_out_281  <= rom_data[281];
			data_out_282  <= rom_data[282];
			data_out_283  <= rom_data[283];
			data_out_284  <= rom_data[284];
			data_out_285  <= rom_data[285];
			data_out_286  <= rom_data[286];
			data_out_287  <= rom_data[287];
			data_out_288  <= rom_data[288];
			data_out_289  <= rom_data[289];
			data_out_290  <= rom_data[290];
			data_out_291  <= rom_data[291];
			data_out_292  <= rom_data[292];
			data_out_293  <= rom_data[293];
			data_out_294  <= rom_data[294];
			data_out_295  <= rom_data[295];
			data_out_296  <= rom_data[296];
			data_out_297  <= rom_data[297];
			data_out_298  <= rom_data[298];
			data_out_299  <= rom_data[299];
			data_out_300  <= rom_data[300];
			data_out_301  <= rom_data[301];
			data_out_302  <= rom_data[302];
			data_out_303  <= rom_data[303];
			data_out_304  <= rom_data[304];
			data_out_305  <= rom_data[305];
			data_out_306  <= rom_data[306];
			data_out_307  <= rom_data[307];
			data_out_308  <= rom_data[308];
			data_out_309  <= rom_data[309];
			data_out_310  <= rom_data[310];
			data_out_311  <= rom_data[311];
			data_out_312  <= rom_data[312];
			data_out_313  <= rom_data[313];
			data_out_314  <= rom_data[314];
			data_out_315  <= rom_data[315];
			data_out_316  <= rom_data[316];
			data_out_317  <= rom_data[317];
			data_out_318  <= rom_data[318];
			data_out_319  <= rom_data[319];
			data_out_320  <= rom_data[320];
			data_out_321  <= rom_data[321];
			data_out_322  <= rom_data[322];
			data_out_323  <= rom_data[323];
			data_out_324  <= rom_data[324];
			data_out_325  <= rom_data[325];
			data_out_326  <= rom_data[326];
			data_out_327  <= rom_data[327];
			data_out_328  <= rom_data[328];
			data_out_329  <= rom_data[329];
			data_out_330  <= rom_data[330];
			data_out_331  <= rom_data[331];
			data_out_332  <= rom_data[332];
			data_out_333  <= rom_data[333];
			data_out_334  <= rom_data[334];
			data_out_335  <= rom_data[335];
			data_out_336  <= rom_data[336];
			data_out_337  <= rom_data[337];
			data_out_338  <= rom_data[338];
			data_out_339  <= rom_data[339];
			data_out_340  <= rom_data[340];
			data_out_341  <= rom_data[341];
			data_out_342  <= rom_data[342];
			data_out_343  <= rom_data[343];
			data_out_344  <= rom_data[344];
			data_out_345  <= rom_data[345];
			data_out_346  <= rom_data[346];
			data_out_347  <= rom_data[347];
			data_out_348  <= rom_data[348];
			data_out_349  <= rom_data[349];
			data_out_350  <= rom_data[350];
			data_out_351  <= rom_data[351];
			data_out_352  <= rom_data[352];
			data_out_353  <= rom_data[353];
			data_out_354  <= rom_data[354];
			data_out_355  <= rom_data[355];
			data_out_356  <= rom_data[356];
			data_out_357  <= rom_data[357];
			data_out_358  <= rom_data[358];
			data_out_359  <= rom_data[359];
			data_out_360  <= rom_data[360];
			data_out_361  <= rom_data[361];
			data_out_362  <= rom_data[362];
			data_out_363  <= rom_data[363];
			data_out_364  <= rom_data[364];
			data_out_365  <= rom_data[365];
			data_out_366  <= rom_data[366];
			data_out_367  <= rom_data[367];
			data_out_368  <= rom_data[368];
			data_out_369  <= rom_data[369];
			data_out_370  <= rom_data[370];
			data_out_371  <= rom_data[371];
			data_out_372  <= rom_data[372];
			data_out_373  <= rom_data[373];
			data_out_374  <= rom_data[374];
			data_out_375  <= rom_data[375];
			data_out_376  <= rom_data[376];
			data_out_377  <= rom_data[377];
			data_out_378  <= rom_data[378];
			data_out_379  <= rom_data[379];
			data_out_380  <= rom_data[380];
			data_out_381  <= rom_data[381];
			data_out_382  <= rom_data[382];
			data_out_383  <= rom_data[383];
			data_out_384  <= rom_data[384];
			data_out_385  <= rom_data[385];
			data_out_386  <= rom_data[386];
			data_out_387  <= rom_data[387];
			data_out_388  <= rom_data[388];
			data_out_389  <= rom_data[389];
			data_out_390  <= rom_data[390];
			data_out_391  <= rom_data[391];
			data_out_392  <= rom_data[392];
			data_out_393  <= rom_data[393];
			data_out_394  <= rom_data[394];
			data_out_395  <= rom_data[395];
			data_out_396  <= rom_data[396];
			data_out_397  <= rom_data[397];
			data_out_398  <= rom_data[398];
			data_out_399  <= rom_data[399];
			data_out_400  <= rom_data[400];
			data_out_401  <= rom_data[401];
			data_out_402  <= rom_data[402];
			data_out_403  <= rom_data[403];
			data_out_404  <= rom_data[404];
			data_out_405  <= rom_data[405];
			data_out_406  <= rom_data[406];
			data_out_407  <= rom_data[407];
			data_out_408  <= rom_data[408];
			data_out_409  <= rom_data[409];
			data_out_410  <= rom_data[410];
			data_out_411  <= rom_data[411];
			data_out_412  <= rom_data[412];
			data_out_413  <= rom_data[413];
			data_out_414  <= rom_data[414];
			data_out_415  <= rom_data[415];
			data_out_416  <= rom_data[416];
			data_out_417  <= rom_data[417];
			data_out_418  <= rom_data[418];
			data_out_419  <= rom_data[419];
			data_out_420  <= rom_data[420];
			data_out_421  <= rom_data[421];
			data_out_422  <= rom_data[422];
			data_out_423  <= rom_data[423];
			data_out_424  <= rom_data[424];
			data_out_425  <= rom_data[425];
			data_out_426  <= rom_data[426];
			data_out_427  <= rom_data[427];
			data_out_428  <= rom_data[428];
			data_out_429  <= rom_data[429];
			data_out_430  <= rom_data[430];
			data_out_431  <= rom_data[431];
			data_out_432  <= rom_data[432];
			data_out_433  <= rom_data[433];
			data_out_434  <= rom_data[434];
			data_out_435  <= rom_data[435];
			data_out_436  <= rom_data[436];
			data_out_437  <= rom_data[437];
			data_out_438  <= rom_data[438];
			data_out_439  <= rom_data[439];
			data_out_440  <= rom_data[440];
			data_out_441  <= rom_data[441];
			data_out_442  <= rom_data[442];
			data_out_443  <= rom_data[443];
			data_out_444  <= rom_data[444];
			data_out_445  <= rom_data[445];
			data_out_446  <= rom_data[446];
			data_out_447  <= rom_data[447];
			data_out_448  <= rom_data[448];
			data_out_449  <= rom_data[449];
			data_out_450  <= rom_data[450];
			data_out_451  <= rom_data[451];
			data_out_452  <= rom_data[452];
			data_out_453  <= rom_data[453];
			data_out_454  <= rom_data[454];
			data_out_455  <= rom_data[455];
			data_out_456  <= rom_data[456];
			data_out_457  <= rom_data[457];
			data_out_458  <= rom_data[458];
			data_out_459  <= rom_data[459];
			data_out_460  <= rom_data[460];
			data_out_461  <= rom_data[461];
			data_out_462  <= rom_data[462];
			data_out_463  <= rom_data[463];
			data_out_464  <= rom_data[464];
			data_out_465  <= rom_data[465];
			data_out_466  <= rom_data[466];
			data_out_467  <= rom_data[467];
			data_out_468  <= rom_data[468];
			data_out_469  <= rom_data[469];
			data_out_470  <= rom_data[470];
			data_out_471  <= rom_data[471];
			data_out_472  <= rom_data[472];
			data_out_473  <= rom_data[473];
			data_out_474  <= rom_data[474];
			data_out_475  <= rom_data[475];
			data_out_476  <= rom_data[476];
			data_out_477  <= rom_data[477];
			data_out_478  <= rom_data[478];
			data_out_479  <= rom_data[479];
			data_out_480  <= rom_data[480];
			data_out_481  <= rom_data[481];
			data_out_482  <= rom_data[482];
			data_out_483  <= rom_data[483];
			data_out_484  <= rom_data[484];
			data_out_485  <= rom_data[485];
			data_out_486  <= rom_data[486];
			data_out_487  <= rom_data[487];
			data_out_488  <= rom_data[488];
			data_out_489  <= rom_data[489];
			data_out_490  <= rom_data[490];
			data_out_491  <= rom_data[491];
			data_out_492  <= rom_data[492];
			data_out_493  <= rom_data[493];
			data_out_494  <= rom_data[494];
			data_out_495  <= rom_data[495];
			data_out_496  <= rom_data[496];
			data_out_497  <= rom_data[497];
			data_out_498  <= rom_data[498];
			data_out_499  <= rom_data[499];
			data_out_500  <= rom_data[500];
			data_out_501  <= rom_data[501];
			data_out_502  <= rom_data[502];
			data_out_503  <= rom_data[503];
			data_out_504  <= rom_data[504];
			data_out_505  <= rom_data[505];
			data_out_506  <= rom_data[506];
			data_out_507  <= rom_data[507];
			data_out_508  <= rom_data[508];
			data_out_509  <= rom_data[509];
			data_out_510  <= rom_data[510];
			data_out_511  <= rom_data[511];
			data_out_512  <= rom_data[512];
			data_out_513  <= rom_data[513];
			data_out_514  <= rom_data[514];
			data_out_515  <= rom_data[515];
			data_out_516  <= rom_data[516];
			data_out_517  <= rom_data[517];
			data_out_518  <= rom_data[518];
			data_out_519  <= rom_data[519];
			data_out_520  <= rom_data[520];
			data_out_521  <= rom_data[521];
			data_out_522  <= rom_data[522];
			data_out_523  <= rom_data[523];
			data_out_524  <= rom_data[524];
			data_out_525  <= rom_data[525];
			data_out_526  <= rom_data[526];
			data_out_527  <= rom_data[527];
			data_out_528  <= rom_data[528];
			data_out_529  <= rom_data[529];
			data_out_530  <= rom_data[530];
			data_out_531  <= rom_data[531];
			data_out_532  <= rom_data[532];
			data_out_533  <= rom_data[533];
			data_out_534  <= rom_data[534];
			data_out_535  <= rom_data[535];
			data_out_536  <= rom_data[536];
			data_out_537  <= rom_data[537];
			data_out_538  <= rom_data[538];
			data_out_539  <= rom_data[539];
			data_out_540  <= rom_data[540];
			data_out_541  <= rom_data[541];
			data_out_542  <= rom_data[542];
			data_out_543  <= rom_data[543];
			data_out_544  <= rom_data[544];
			data_out_545  <= rom_data[545];
			data_out_546  <= rom_data[546];
			data_out_547  <= rom_data[547];
			data_out_548  <= rom_data[548];
			data_out_549  <= rom_data[549];
			data_out_550  <= rom_data[550];
			data_out_551  <= rom_data[551];
			data_out_552  <= rom_data[552];
			data_out_553  <= rom_data[553];
			data_out_554  <= rom_data[554];
			data_out_555  <= rom_data[555];
			data_out_556  <= rom_data[556];
			data_out_557  <= rom_data[557];
			data_out_558  <= rom_data[558];
			data_out_559  <= rom_data[559];
			data_out_560  <= rom_data[560];
			data_out_561  <= rom_data[561];
			data_out_562  <= rom_data[562];
			data_out_563  <= rom_data[563];
			data_out_564  <= rom_data[564];
			data_out_565  <= rom_data[565];
			data_out_566  <= rom_data[566];
			data_out_567  <= rom_data[567];
			data_out_568  <= rom_data[568];
			data_out_569  <= rom_data[569];
			data_out_570  <= rom_data[570];
			data_out_571  <= rom_data[571];
			data_out_572  <= rom_data[572];
			data_out_573  <= rom_data[573];
			data_out_574  <= rom_data[574];
			data_out_575  <= rom_data[575];
			data_out_576  <= rom_data[576];
			data_out_577  <= rom_data[577];
			data_out_578  <= rom_data[578];
			data_out_579  <= rom_data[579];
			data_out_580  <= rom_data[580];
			data_out_581  <= rom_data[581];
			data_out_582  <= rom_data[582];
			data_out_583  <= rom_data[583];
			data_out_584  <= rom_data[584];
			data_out_585  <= rom_data[585];
			data_out_586  <= rom_data[586];
			data_out_587  <= rom_data[587];
			data_out_588  <= rom_data[588];
			data_out_589  <= rom_data[589];
			data_out_590  <= rom_data[590];
			data_out_591  <= rom_data[591];
			data_out_592  <= rom_data[592];
			data_out_593  <= rom_data[593];
			data_out_594  <= rom_data[594];
			data_out_595  <= rom_data[595];
			data_out_596  <= rom_data[596];
			data_out_597  <= rom_data[597];
			data_out_598  <= rom_data[598];
			data_out_599  <= rom_data[599];
			data_out_600  <= rom_data[600];
			data_out_601  <= rom_data[601];
			data_out_602  <= rom_data[602];
			data_out_603  <= rom_data[603];
			data_out_604  <= rom_data[604];
			data_out_605  <= rom_data[605];
			data_out_606  <= rom_data[606];
			data_out_607  <= rom_data[607];
			data_out_608  <= rom_data[608];
			data_out_609  <= rom_data[609];
			data_out_610  <= rom_data[610];
			data_out_611  <= rom_data[611];
			data_out_612  <= rom_data[612];
			data_out_613  <= rom_data[613];
			data_out_614  <= rom_data[614];
			data_out_615  <= rom_data[615];
			data_out_616  <= rom_data[616];
			data_out_617  <= rom_data[617];
			data_out_618  <= rom_data[618];
			data_out_619  <= rom_data[619];
			data_out_620  <= rom_data[620];
			data_out_621  <= rom_data[621];
			data_out_622  <= rom_data[622];
			data_out_623  <= rom_data[623];
			data_out_624  <= rom_data[624];
			data_out_625  <= rom_data[625];
			data_out_626  <= rom_data[626];
			data_out_627  <= rom_data[627];
			data_out_628  <= rom_data[628];
			data_out_629  <= rom_data[629];
			data_out_630  <= rom_data[630];
			data_out_631  <= rom_data[631];
			data_out_632  <= rom_data[632];
			data_out_633  <= rom_data[633];
			data_out_634  <= rom_data[634];
			data_out_635  <= rom_data[635];
			data_out_636  <= rom_data[636];
			data_out_637  <= rom_data[637];
			data_out_638  <= rom_data[638];
			data_out_639  <= rom_data[639];
			data_out_640  <= rom_data[640];
			data_out_641  <= rom_data[641];
			data_out_642  <= rom_data[642];
			data_out_643  <= rom_data[643];
			data_out_644  <= rom_data[644];
			data_out_645  <= rom_data[645];
			data_out_646  <= rom_data[646];
			data_out_647  <= rom_data[647];
			data_out_648  <= rom_data[648];
			data_out_649  <= rom_data[649];
			data_out_650  <= rom_data[650];
			data_out_651  <= rom_data[651];
			data_out_652  <= rom_data[652];
			data_out_653  <= rom_data[653];
			data_out_654  <= rom_data[654];
			data_out_655  <= rom_data[655];
			data_out_656  <= rom_data[656];
			data_out_657  <= rom_data[657];
			data_out_658  <= rom_data[658];
			data_out_659  <= rom_data[659];
			data_out_660  <= rom_data[660];
			data_out_661  <= rom_data[661];
			data_out_662  <= rom_data[662];
			data_out_663  <= rom_data[663];
			data_out_664  <= rom_data[664];
			data_out_665  <= rom_data[665];
			data_out_666  <= rom_data[666];
			data_out_667  <= rom_data[667];
			data_out_668  <= rom_data[668];
			data_out_669  <= rom_data[669];
			data_out_670  <= rom_data[670];
			data_out_671  <= rom_data[671];
			data_out_672  <= rom_data[672];
			data_out_673  <= rom_data[673];
			data_out_674  <= rom_data[674];
			data_out_675  <= rom_data[675];
			data_out_676  <= rom_data[676];
			data_out_677  <= rom_data[677];
			data_out_678  <= rom_data[678];
			data_out_679  <= rom_data[679];
			data_out_680  <= rom_data[680];
			data_out_681  <= rom_data[681];
			data_out_682  <= rom_data[682];
			data_out_683  <= rom_data[683];
			data_out_684  <= rom_data[684];
			data_out_685  <= rom_data[685];
			data_out_686  <= rom_data[686];
			data_out_687  <= rom_data[687];
			data_out_688  <= rom_data[688];
			data_out_689  <= rom_data[689];
			data_out_690  <= rom_data[690];
			data_out_691  <= rom_data[691];
			data_out_692  <= rom_data[692];
			data_out_693  <= rom_data[693];
			data_out_694  <= rom_data[694];
			data_out_695  <= rom_data[695];
			data_out_696  <= rom_data[696];
			data_out_697  <= rom_data[697];
			data_out_698  <= rom_data[698];
			data_out_699  <= rom_data[699];
			data_out_700  <= rom_data[700];
			data_out_701  <= rom_data[701];
			data_out_702  <= rom_data[702];
			data_out_703  <= rom_data[703];
			data_out_704  <= rom_data[704];
			data_out_705  <= rom_data[705];
			data_out_706  <= rom_data[706];
			data_out_707  <= rom_data[707];
			data_out_708  <= rom_data[708];
			data_out_709  <= rom_data[709];
			data_out_710  <= rom_data[710];
			data_out_711  <= rom_data[711];
			data_out_712  <= rom_data[712];
			data_out_713  <= rom_data[713];
			data_out_714  <= rom_data[714];
			data_out_715  <= rom_data[715];
			data_out_716  <= rom_data[716];
			data_out_717  <= rom_data[717];
			data_out_718  <= rom_data[718];
			data_out_719  <= rom_data[719];
			data_out_720  <= rom_data[720];
			data_out_721  <= rom_data[721];
			data_out_722  <= rom_data[722];
			data_out_723  <= rom_data[723];
			data_out_724  <= rom_data[724];
			data_out_725  <= rom_data[725];
			data_out_726  <= rom_data[726];
			data_out_727  <= rom_data[727];
			data_out_728  <= rom_data[728];
			data_out_729  <= rom_data[729];
			data_out_730  <= rom_data[730];
			data_out_731  <= rom_data[731];
			data_out_732  <= rom_data[732];
			data_out_733  <= rom_data[733];
			data_out_734  <= rom_data[734];
			data_out_735  <= rom_data[735];
			data_out_736  <= rom_data[736];
			data_out_737  <= rom_data[737];
			data_out_738  <= rom_data[738];
			data_out_739  <= rom_data[739];


        end
    end
endmodule
