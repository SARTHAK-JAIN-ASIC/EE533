module tb_NPU_pipeline_top;

   reg clk;
   reg reset;
   reg [63:0] data_in;
   reg valid_in;

   NPU_pipeline_top uut(
	.clk(clk),
	.reset(reset),
	.data_in(data_in),
	.valid_in(valid_in)
	// .data_in(64'b0011110000111100001011000000110000000110000000100010011000111100)
   );
   
  /*  initial
   begin
	  reset      = 0;
	  clk        = 0;
	  #80; reset = ~reset;
	  #80; reset = ~reset;
		#10000;
      $finish;
	end */

	always
	begin
		#10 clk = ~clk;
	end
	
	initial begin
	  reset      = 0;
	  clk        = 0;
	  data_in    = 0;
	  valid_in   = 0;
	  #80; reset = ~reset;
	  #80; reset = ~reset;
	  // #40;
    
	// Actual: 1
	valid_in   = 1;
	data_in = 64'b0001100000111000011111000100100000011000000110000001100000011000;
    #1300;  // Wait 65 clocks
	
	// Actual: 2
    data_in = 64'b0011100000111000000011000000100000001000001110000011110000110000;
    #1300;  // Wait 65 clocks
	
	 // Actual: 0
    data_in = 64'b0001100000111100001001000000000000000000001001000011110000011000;
    #1300;  // Wait 65 clocks
	
	// Actual: 2
    data_in = 64'b0001100001111000011010000000110000001000000010000001111000011111;
    #1300;  // Wait 65 clocks
	
	// valid_in = 0;
	
	// Actual: 4
    data_in = 64'b0000100000011100000101000010110000111100000111000000100000001000;
    #1300;  // Wait 65 clocks
	
	// valid_in = 0;
	
	// Actual: 3
	data_in = 64'b0011110000111100001011000000110000000110000000100010011000111100;
    #1300;  // Wait 65 clocks
	
	// valid_in = 0;
	
	// Actual: 5
    data_in = 64'b0000111000111100001000000011100000001100000011000011100000110000;
    #1300;  // Wait 65 clocks
	
	// valid_in = 0;
	
	 // Actual: 7
    data_in = 64'b0001111000111110001000100010010000001000000010000001100000010000;
    #1300;  // Wait 65 clocks
	
	// Actual: 2
    data_in = 64'b0011000000111000011010000000100000011000000100000011111000110000;
    #1300;  // Wait 65 clocks
	
	// Actual: 1
    data_in = 64'b0000010000001110000111000011110000001100000011000000110000000100;
    #1300;  // Wait 65 clocks  

 






 
   /*  // Actual: 6
	data_in = 64'b0001000000110000001000000010000000100000001111100011011000011100;
    #1300;  // Wait 65 clocks
	
	// Actual: 3
    data_in = 64'b0011100000101000000001000001100000011100000001000110010000011100;
    #1300;  // Wait 65 clocks
	
	 // Actual: 4
    data_in = 64'b0001100000110000001000000010010000111100000011000000100000011000;
    #1300;  // Wait 65 clocks
	
	// Actual: 0
    data_in = 64'b0011100000111000001001000010010000100000001000000010010000011100;
    #1300;  // Wait 65 clocks
	
	// Actual: 2
    data_in = 64'b0011100000111000001111000000100000001000000110000011101000111111;
    #1300;  // Wait 65 clocks
	
	// Actual: 2
	data_in = 64'b0001100000011100000001000000010000001100000011000001111100011100;
    #1300;  // Wait 65 clocks
	
	// Actual: 2
    data_in = 64'b0011100000101000000010000000100000011000000100000011110000111000;
    #1300;  // Wait 65 clocks
	
	 // Actual: 7
    data_in = 64'b0001110000111100001010000000100000011110000110000001000000010000;
    #1300;  // Wait 65 clocks
	
	// Actual: 3
    data_in = 64'b0011100000101100000010000001100000001100000001000000010000111100;
    #1300;  // Wait 65 clocks
	
	// Actual: 3
    data_in = 64'b0001100000101100000010000001100000000100000001000010010000111000;
    #1300;  // Wait 65 clocks   */
 
 
 
	
	
	
	
	
	
	


	
	#1000 //Run for another 1000 ns

    // End the simulation
    $finish;
  end


endmodule
